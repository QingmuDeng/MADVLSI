magic
tech sky130A
timestamp 1612836255
<< locali >>
rect -120 -40 -100 -20
rect 270 -40 290 -20
<< metal1 >>
rect -120 155 -100 245
rect -120 0 -100 90
use inverter  inverter_1
timestamp 1612836176
transform 1 0 615 0 1 140
box -530 -200 -325 130
use inverter  inverter_0
timestamp 1612836176
transform 1 0 410 0 1 140
box -530 -200 -325 130
<< labels >>
rlabel locali -120 -30 -120 -30 7 A
rlabel locali 290 -30 290 -30 3 Y
rlabel metal1 -120 45 -120 45 7 VN
rlabel metal1 -120 195 -120 195 7 VP
<< end >>
