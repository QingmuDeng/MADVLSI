magic
tech sky130A
timestamp 1612836176
<< nwell >>
rect -530 -10 -325 130
<< nmos >>
rect -410 -145 -395 -45
<< pmos >>
rect -410 10 -395 110
<< ndiff >>
rect -460 -60 -410 -45
rect -460 -130 -445 -60
rect -425 -130 -410 -60
rect -460 -145 -410 -130
rect -395 -60 -345 -45
rect -395 -130 -380 -60
rect -360 -130 -345 -60
rect -395 -145 -345 -130
<< pdiff >>
rect -460 95 -410 110
rect -460 25 -445 95
rect -425 25 -410 95
rect -460 10 -410 25
rect -395 95 -345 110
rect -395 25 -380 95
rect -360 25 -345 95
rect -395 10 -345 25
<< ndiffc >>
rect -445 -130 -425 -60
rect -380 -130 -360 -60
<< pdiffc >>
rect -445 25 -425 95
rect -380 25 -360 95
<< psubdiff >>
rect -510 -60 -460 -45
rect -510 -130 -495 -60
rect -475 -130 -460 -60
rect -510 -145 -460 -130
<< nsubdiff >>
rect -510 95 -460 110
rect -510 25 -495 95
rect -475 25 -460 95
rect -510 10 -460 25
<< psubdiffcont >>
rect -495 -130 -475 -60
<< nsubdiffcont >>
rect -495 25 -475 95
<< poly >>
rect -410 110 -395 125
rect -410 -45 -395 10
rect -410 -160 -395 -145
rect -435 -170 -395 -160
rect -435 -190 -425 -170
rect -405 -190 -395 -170
rect -435 -200 -395 -190
<< polycont >>
rect -425 -190 -405 -170
<< locali >>
rect -505 95 -415 105
rect -505 25 -495 95
rect -475 25 -445 95
rect -425 25 -415 95
rect -505 15 -415 25
rect -390 95 -350 105
rect -390 25 -380 95
rect -360 25 -350 95
rect -390 15 -350 25
rect -370 -50 -350 15
rect -505 -60 -415 -50
rect -505 -130 -495 -60
rect -475 -130 -445 -60
rect -425 -130 -415 -60
rect -505 -140 -415 -130
rect -390 -60 -350 -50
rect -390 -130 -380 -60
rect -360 -130 -350 -60
rect -390 -140 -350 -130
rect -370 -160 -350 -140
rect -530 -170 -395 -160
rect -530 -180 -425 -170
rect -435 -190 -425 -180
rect -405 -190 -395 -170
rect -370 -180 -325 -160
rect -435 -200 -395 -190
<< viali >>
rect -495 25 -475 95
rect -445 25 -425 95
rect -495 -130 -475 -60
rect -445 -130 -425 -60
<< metal1 >>
rect -530 95 -325 105
rect -530 25 -495 95
rect -475 25 -445 95
rect -425 25 -325 95
rect -530 15 -325 25
rect -530 -60 -325 -50
rect -530 -130 -495 -60
rect -475 -130 -445 -60
rect -425 -130 -325 -60
rect -530 -140 -325 -130
<< labels >>
rlabel space -510 -160 -345 -30 1 :
rlabel locali -530 -170 -530 -170 7 A
port 1 w
rlabel locali -325 -170 -325 -170 3 Y
port 2 e
rlabel metal1 -530 -96 -530 -95 7 VN
port 4 w
rlabel metal1 -530 60 -530 60 7 VP
port 3 w
<< end >>
