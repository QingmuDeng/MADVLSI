magic
tech sky130A
timestamp 1612889628
<< nwell >>
rect -145 135 125 275
<< nmos >>
rect 0 0 15 100
rect 40 0 55 100
<< pmos >>
rect -25 155 -10 255
rect 40 155 55 255
<< ndiff >>
rect -50 85 0 100
rect -50 15 -35 85
rect -15 15 0 85
rect -50 0 0 15
rect 15 0 40 100
rect 55 85 105 100
rect 55 15 70 85
rect 90 15 105 85
rect 55 0 105 15
<< pdiff >>
rect -75 240 -25 255
rect -75 170 -60 240
rect -40 170 -25 240
rect -75 155 -25 170
rect -10 240 40 255
rect -10 170 5 240
rect 25 170 40 240
rect -10 155 40 170
rect 55 240 105 255
rect 55 170 70 240
rect 90 170 105 240
rect 55 155 105 170
<< ndiffc >>
rect -35 15 -15 85
rect 70 15 90 85
<< pdiffc >>
rect -60 170 -40 240
rect 5 170 25 240
rect 70 170 90 240
<< psubdiff >>
rect -125 85 -50 100
rect -125 15 -110 85
rect -90 15 -50 85
rect -125 0 -50 15
<< nsubdiff >>
rect -125 240 -75 255
rect -125 170 -110 240
rect -90 170 -75 240
rect -125 155 -75 170
<< psubdiffcont >>
rect -110 15 -90 85
<< nsubdiffcont >>
rect -110 170 -90 240
<< poly >>
rect 15 300 55 310
rect 15 280 25 300
rect 45 280 55 300
rect 15 270 55 280
rect -25 255 -10 270
rect 40 255 55 270
rect -25 135 -10 155
rect -25 120 15 135
rect 0 100 15 120
rect 40 100 55 155
rect 0 -15 15 0
rect 40 -15 55 0
rect -25 -25 15 -15
rect -25 -45 -15 -25
rect 5 -45 15 -25
rect -25 -55 15 -45
<< polycont >>
rect 25 280 45 300
rect -15 -45 5 -25
<< locali >>
rect 15 300 55 310
rect 15 290 25 300
rect -145 280 25 290
rect 45 280 55 300
rect -145 270 55 280
rect -120 240 -30 250
rect -120 170 -110 240
rect -90 170 -60 240
rect -40 170 -30 240
rect -120 160 -30 170
rect -5 240 35 250
rect -5 170 5 240
rect 25 170 35 240
rect -5 160 35 170
rect 60 240 100 250
rect 60 170 70 240
rect 90 170 100 240
rect 60 160 100 170
rect 15 135 35 160
rect 15 115 100 135
rect 80 95 100 115
rect -120 85 -5 95
rect -120 15 -110 85
rect -90 15 -35 85
rect -15 15 -5 85
rect -120 5 -5 15
rect 60 85 100 95
rect 60 15 70 85
rect 90 15 100 85
rect 60 5 100 15
rect 80 -15 100 5
rect -145 -25 15 -15
rect -145 -35 -15 -25
rect -25 -45 -15 -35
rect 5 -45 15 -25
rect 80 -35 125 -15
rect -25 -55 15 -45
<< viali >>
rect -110 170 -90 240
rect -60 170 -40 240
rect 70 170 90 240
rect -110 15 -90 85
rect -35 15 -15 85
<< metal1 >>
rect -145 240 125 250
rect -145 170 -110 240
rect -90 170 -60 240
rect -40 170 70 240
rect 90 170 125 240
rect -145 160 125 170
rect -145 85 125 95
rect -145 15 -110 85
rect -90 15 -35 85
rect -15 15 125 85
rect -145 5 125 15
<< labels >>
rlabel locali -145 -25 -145 -25 7 A
port 1 w
rlabel locali 125 -25 125 -25 3 Y
port 3 e
rlabel metal1 -145 205 -145 205 7 VP
port 4 w
rlabel locali -145 280 -145 280 7 B
port 2 w
rlabel metal1 -145 50 -145 50 7 VN
port 5 w
<< end >>
