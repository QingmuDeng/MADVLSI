magic
tech sky130A
timestamp 1615258683
<< nmos >>
rect -400 3365 -350 3965
rect -300 3365 -250 3965
rect -200 3365 -150 3965
rect -100 3365 -50 3965
rect 0 3365 50 3965
rect 100 3365 150 3965
rect 200 3365 250 3965
rect 300 3365 350 3965
rect 400 3365 450 3965
rect 500 3365 550 3965
rect -400 2065 -350 3265
rect -300 2065 -250 3265
rect -200 2065 -150 3265
rect -100 2065 -50 3265
rect 0 2065 50 3265
rect 100 2065 150 3265
rect 200 2065 250 3265
rect 300 2065 350 3265
rect 400 2065 450 3265
rect 500 2065 550 3265
rect -395 1315 -345 1915
rect -295 1315 -245 1915
rect -195 1315 -145 1915
rect -95 1315 -45 1915
rect 5 1315 55 1915
rect 105 1315 155 1915
rect 205 1315 255 1915
rect 305 1315 355 1915
rect 405 1315 455 1915
rect 505 1315 555 1915
rect -395 315 -345 915
rect -295 315 -245 915
rect -195 315 -145 915
rect -95 315 -45 915
rect 5 315 55 915
rect 105 315 155 915
rect 205 315 255 915
rect 305 315 355 915
rect 405 315 455 915
rect 505 315 555 915
<< ndiff >>
rect -450 3950 -400 3965
rect -450 3380 -435 3950
rect -415 3380 -400 3950
rect -450 3365 -400 3380
rect -350 3950 -300 3965
rect -350 3380 -335 3950
rect -315 3380 -300 3950
rect -350 3365 -300 3380
rect -250 3950 -200 3965
rect -250 3380 -235 3950
rect -215 3380 -200 3950
rect -250 3365 -200 3380
rect -150 3950 -100 3965
rect -150 3380 -135 3950
rect -115 3380 -100 3950
rect -150 3365 -100 3380
rect -50 3950 0 3965
rect -50 3380 -35 3950
rect -15 3380 0 3950
rect -50 3365 0 3380
rect 50 3950 100 3965
rect 50 3380 65 3950
rect 85 3380 100 3950
rect 50 3365 100 3380
rect 150 3950 200 3965
rect 150 3380 165 3950
rect 185 3380 200 3950
rect 150 3365 200 3380
rect 250 3950 300 3965
rect 250 3380 265 3950
rect 285 3380 300 3950
rect 250 3365 300 3380
rect 350 3950 400 3965
rect 350 3380 365 3950
rect 385 3380 400 3950
rect 350 3365 400 3380
rect 450 3950 500 3965
rect 450 3380 465 3950
rect 485 3380 500 3950
rect 450 3365 500 3380
rect 550 3950 600 3965
rect 550 3380 565 3950
rect 585 3380 600 3950
rect 550 3365 600 3380
rect -450 3245 -400 3265
rect -450 2080 -435 3245
rect -415 2080 -400 3245
rect -450 2065 -400 2080
rect -350 3245 -300 3265
rect -350 2080 -335 3245
rect -315 2080 -300 3245
rect -350 2065 -300 2080
rect -250 3245 -200 3265
rect -250 2080 -235 3245
rect -215 2080 -200 3245
rect -250 2065 -200 2080
rect -150 3245 -100 3265
rect -150 2080 -135 3245
rect -115 2080 -100 3245
rect -150 2065 -100 2080
rect -50 3245 0 3265
rect -50 2080 -35 3245
rect -15 2080 0 3245
rect -50 2065 0 2080
rect 50 3245 100 3265
rect 50 2080 65 3245
rect 85 2080 100 3245
rect 50 2065 100 2080
rect 150 3245 200 3265
rect 150 2080 165 3245
rect 185 2080 200 3245
rect 150 2065 200 2080
rect 250 3245 300 3265
rect 250 2080 265 3245
rect 285 2080 300 3245
rect 250 2065 300 2080
rect 350 3245 400 3265
rect 350 2080 365 3245
rect 385 2080 400 3245
rect 350 2065 400 2080
rect 450 3245 500 3265
rect 450 2080 465 3245
rect 485 2080 500 3245
rect 450 2065 500 2080
rect 550 3245 600 3265
rect 550 2080 565 3245
rect 585 2080 600 3245
rect 550 2065 600 2080
rect -445 1900 -395 1915
rect -445 1330 -430 1900
rect -410 1330 -395 1900
rect -445 1315 -395 1330
rect -345 1900 -295 1915
rect -345 1330 -330 1900
rect -310 1330 -295 1900
rect -345 1315 -295 1330
rect -245 1900 -195 1915
rect -245 1330 -230 1900
rect -210 1330 -195 1900
rect -245 1315 -195 1330
rect -145 1900 -95 1915
rect -145 1330 -130 1900
rect -110 1330 -95 1900
rect -145 1315 -95 1330
rect -45 1900 5 1915
rect -45 1330 -30 1900
rect -10 1330 5 1900
rect -45 1315 5 1330
rect 55 1900 105 1915
rect 55 1330 70 1900
rect 90 1330 105 1900
rect 55 1315 105 1330
rect 155 1900 205 1915
rect 155 1330 170 1900
rect 190 1330 205 1900
rect 155 1315 205 1330
rect 255 1900 305 1915
rect 255 1330 270 1900
rect 290 1330 305 1900
rect 255 1315 305 1330
rect 355 1900 405 1915
rect 355 1330 370 1900
rect 390 1330 405 1900
rect 355 1315 405 1330
rect 455 1900 505 1915
rect 455 1330 470 1900
rect 490 1330 505 1900
rect 455 1315 505 1330
rect 555 1900 605 1915
rect 555 1330 570 1900
rect 590 1330 605 1900
rect 555 1315 605 1330
rect -445 900 -395 915
rect -445 330 -430 900
rect -410 330 -395 900
rect -445 315 -395 330
rect -345 900 -295 915
rect -345 330 -330 900
rect -310 330 -295 900
rect -345 315 -295 330
rect -245 900 -195 915
rect -245 330 -230 900
rect -210 330 -195 900
rect -245 315 -195 330
rect -145 900 -95 915
rect -145 330 -130 900
rect -110 330 -95 900
rect -145 315 -95 330
rect -45 900 5 915
rect -45 330 -30 900
rect -10 330 5 900
rect -45 315 5 330
rect 55 900 105 915
rect 55 330 70 900
rect 90 330 105 900
rect 55 315 105 330
rect 155 900 205 915
rect 155 330 170 900
rect 190 330 205 900
rect 155 315 205 330
rect 255 900 305 915
rect 255 330 270 900
rect 290 330 305 900
rect 255 315 305 330
rect 355 900 405 915
rect 355 330 370 900
rect 390 330 405 900
rect 355 315 405 330
rect 455 900 505 915
rect 455 330 470 900
rect 490 330 505 900
rect 455 315 505 330
rect 555 900 605 915
rect 555 330 570 900
rect 590 330 605 900
rect 555 315 605 330
<< ndiffc >>
rect -435 3380 -415 3950
rect -335 3380 -315 3950
rect -235 3380 -215 3950
rect -135 3380 -115 3950
rect -35 3380 -15 3950
rect 65 3380 85 3950
rect 165 3380 185 3950
rect 265 3380 285 3950
rect 365 3380 385 3950
rect 465 3380 485 3950
rect 565 3380 585 3950
rect -435 2080 -415 3245
rect -335 2080 -315 3245
rect -235 2080 -215 3245
rect -135 2080 -115 3245
rect -35 2080 -15 3245
rect 65 2080 85 3245
rect 165 2080 185 3245
rect 265 2080 285 3245
rect 365 2080 385 3245
rect 465 2080 485 3245
rect 565 2080 585 3245
rect -430 1330 -410 1900
rect -330 1330 -310 1900
rect -230 1330 -210 1900
rect -130 1330 -110 1900
rect -30 1330 -10 1900
rect 70 1330 90 1900
rect 170 1330 190 1900
rect 270 1330 290 1900
rect 370 1330 390 1900
rect 470 1330 490 1900
rect 570 1330 590 1900
rect -430 330 -410 900
rect -330 330 -310 900
rect -230 330 -210 900
rect -130 330 -110 900
rect -30 330 -10 900
rect 70 330 90 900
rect 170 330 190 900
rect 270 330 290 900
rect 370 330 390 900
rect 470 330 490 900
rect 570 330 590 900
<< poly >>
rect -400 3965 -350 3980
rect -300 3965 -250 3980
rect -200 3965 -150 3980
rect -100 3965 -50 3980
rect 0 3965 50 3980
rect 100 3965 150 3980
rect 200 3965 250 3980
rect 300 3965 350 3980
rect 400 3965 450 3980
rect 500 3965 550 3980
rect -400 3350 -350 3365
rect -300 3350 -250 3365
rect -200 3350 -150 3365
rect -100 3350 -50 3365
rect 0 3350 50 3365
rect 100 3350 150 3365
rect 200 3350 250 3365
rect 300 3350 350 3365
rect 400 3350 450 3365
rect 500 3350 550 3365
rect -400 3265 -350 3280
rect -300 3265 -250 3280
rect -200 3265 -150 3280
rect -100 3265 -50 3280
rect 0 3265 50 3280
rect 100 3265 150 3280
rect 200 3265 250 3280
rect 300 3265 350 3280
rect 400 3265 450 3280
rect 500 3265 550 3280
rect -400 2050 -350 2065
rect -300 2050 -250 2065
rect -200 2050 -150 2065
rect -100 2050 -50 2065
rect 0 2050 50 2065
rect 100 2050 150 2065
rect 200 2050 250 2065
rect 300 2050 350 2065
rect 400 2050 450 2065
rect 500 2050 550 2065
rect -395 1915 -345 1930
rect -295 1915 -245 1930
rect -195 1915 -145 1930
rect -95 1915 -45 1930
rect 5 1915 55 1930
rect 105 1915 155 1930
rect 205 1915 255 1930
rect 305 1915 355 1930
rect 405 1915 455 1930
rect 505 1915 555 1930
rect -395 1300 -345 1315
rect -295 1300 -245 1315
rect -195 1300 -145 1315
rect -95 1300 -45 1315
rect 5 1300 55 1315
rect 105 1300 155 1315
rect 205 1300 255 1315
rect 305 1300 355 1315
rect 405 1300 455 1315
rect 505 1300 555 1315
rect -395 915 -345 930
rect -295 915 -245 930
rect -195 915 -145 930
rect -95 915 -45 930
rect 5 915 55 930
rect 105 915 155 930
rect 205 915 255 930
rect 305 915 355 930
rect 405 915 455 930
rect 505 915 555 930
rect -395 300 -345 315
rect -295 300 -245 315
rect -195 300 -145 315
rect -95 300 -45 315
rect 5 300 55 315
rect 105 300 155 315
rect 205 300 255 315
rect 305 300 355 315
rect 405 300 455 315
rect 505 300 555 315
<< locali >>
rect -445 3950 -405 3960
rect -445 3380 -435 3950
rect -415 3380 -405 3950
rect -445 3370 -405 3380
rect -345 3950 -305 3960
rect -345 3380 -335 3950
rect -315 3380 -305 3950
rect -345 3370 -305 3380
rect -245 3950 -205 3960
rect -245 3380 -235 3950
rect -215 3380 -205 3950
rect -245 3370 -205 3380
rect -145 3950 -105 3960
rect -145 3380 -135 3950
rect -115 3380 -105 3950
rect -145 3370 -105 3380
rect -45 3950 -5 3960
rect -45 3380 -35 3950
rect -15 3380 -5 3950
rect -45 3370 -5 3380
rect 55 3950 95 3960
rect 55 3380 65 3950
rect 85 3380 95 3950
rect 55 3370 95 3380
rect 155 3950 195 3960
rect 155 3380 165 3950
rect 185 3380 195 3950
rect 155 3370 195 3380
rect 255 3950 295 3960
rect 255 3380 265 3950
rect 285 3380 295 3950
rect 255 3370 295 3380
rect 355 3950 395 3960
rect 355 3380 365 3950
rect 385 3380 395 3950
rect 355 3370 395 3380
rect 455 3950 495 3960
rect 455 3380 465 3950
rect 485 3380 495 3950
rect 455 3370 495 3380
rect 555 3950 595 3960
rect 555 3380 565 3950
rect 585 3380 595 3950
rect 555 3370 595 3380
rect -445 3245 -405 3255
rect -445 2080 -435 3245
rect -415 2080 -405 3245
rect -445 2070 -405 2080
rect -345 3245 -305 3255
rect -345 2080 -335 3245
rect -315 2080 -305 3245
rect -345 2070 -305 2080
rect -245 3245 -205 3255
rect -245 2080 -235 3245
rect -215 2080 -205 3245
rect -245 2070 -205 2080
rect -145 3245 -105 3255
rect -145 2080 -135 3245
rect -115 2080 -105 3245
rect -145 2070 -105 2080
rect -45 3245 -5 3255
rect -45 2080 -35 3245
rect -15 2080 -5 3245
rect -45 2070 -5 2080
rect 55 3245 95 3255
rect 55 2080 65 3245
rect 85 2080 95 3245
rect 55 2070 95 2080
rect 155 3245 195 3255
rect 155 2080 165 3245
rect 185 2080 195 3245
rect 155 2070 195 2080
rect 255 3245 295 3255
rect 255 2080 265 3245
rect 285 2080 295 3245
rect 255 2070 295 2080
rect 355 3245 395 3255
rect 355 2080 365 3245
rect 385 2080 395 3245
rect 355 2070 395 2080
rect 455 3245 495 3255
rect 455 2080 465 3245
rect 485 2080 495 3245
rect 455 2070 495 2080
rect 555 3245 595 3255
rect 555 2080 565 3245
rect 585 2080 595 3245
rect 555 2070 595 2080
rect -440 1900 -400 1910
rect -440 1330 -430 1900
rect -410 1330 -400 1900
rect -440 1320 -400 1330
rect -340 1900 -300 1910
rect -340 1330 -330 1900
rect -310 1330 -300 1900
rect -340 1320 -300 1330
rect -240 1900 -200 1910
rect -240 1330 -230 1900
rect -210 1330 -200 1900
rect -240 1320 -200 1330
rect -140 1900 -100 1910
rect -140 1330 -130 1900
rect -110 1330 -100 1900
rect -140 1320 -100 1330
rect -40 1900 0 1910
rect -40 1330 -30 1900
rect -10 1330 0 1900
rect -40 1320 0 1330
rect 60 1900 100 1910
rect 60 1330 70 1900
rect 90 1330 100 1900
rect 60 1320 100 1330
rect 160 1900 200 1910
rect 160 1330 170 1900
rect 190 1330 200 1900
rect 160 1320 200 1330
rect 260 1900 300 1910
rect 260 1330 270 1900
rect 290 1330 300 1900
rect 260 1320 300 1330
rect 360 1900 400 1910
rect 360 1330 370 1900
rect 390 1330 400 1900
rect 360 1320 400 1330
rect 460 1900 500 1910
rect 460 1330 470 1900
rect 490 1330 500 1900
rect 460 1320 500 1330
rect 560 1900 600 1910
rect 560 1330 570 1900
rect 590 1330 600 1900
rect 560 1320 600 1330
rect -440 900 -400 910
rect -440 330 -430 900
rect -410 330 -400 900
rect -440 320 -400 330
rect -340 900 -300 910
rect -340 330 -330 900
rect -310 330 -300 900
rect -340 320 -300 330
rect -240 900 -200 910
rect -240 330 -230 900
rect -210 330 -200 900
rect -240 320 -200 330
rect -140 900 -100 910
rect -140 330 -130 900
rect -110 330 -100 900
rect -140 320 -100 330
rect -40 900 0 910
rect -40 330 -30 900
rect -10 330 0 900
rect -40 320 0 330
rect 60 900 100 910
rect 60 330 70 900
rect 90 330 100 900
rect 60 320 100 330
rect 160 900 200 910
rect 160 330 170 900
rect 190 330 200 900
rect 160 320 200 330
rect 260 900 300 910
rect 260 330 270 900
rect 290 330 300 900
rect 260 320 300 330
rect 360 900 400 910
rect 360 330 370 900
rect 390 330 400 900
rect 360 320 400 330
rect 460 900 500 910
rect 460 330 470 900
rect 490 330 500 900
rect 460 320 500 330
rect 560 900 600 910
rect 560 330 570 900
rect 590 330 600 900
rect 560 320 600 330
<< end >>
