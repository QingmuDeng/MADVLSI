magic
tech sky130A
timestamp 1615435668
<< nwell >>
rect -2415 1290 580 1930
<< nmos >>
rect -2295 380 -2245 980
rect -2195 380 -2145 980
rect -2095 380 -2045 980
rect -1995 380 -1945 980
rect -1895 380 -1845 980
rect -1795 380 -1745 980
rect -1595 380 -1545 980
rect -1495 380 -1445 980
rect -1395 380 -1345 980
rect -1295 380 -1245 980
rect -1195 380 -1145 980
rect -1095 380 -1045 980
rect -995 380 -945 980
rect -895 380 -845 980
rect -795 380 -745 980
rect -695 380 -645 980
rect -495 380 -445 980
rect -395 380 -345 980
rect -295 380 -245 980
rect -195 380 -145 980
rect -95 380 -45 980
rect 5 380 55 980
rect 105 380 155 980
rect 205 380 255 980
rect 305 380 355 980
rect 405 380 455 980
<< pmos >>
rect -2295 1310 -2245 1910
rect -2195 1310 -2145 1910
rect -2095 1310 -2045 1910
rect -1995 1310 -1945 1910
rect -1895 1310 -1845 1910
rect -1795 1310 -1745 1910
rect -1595 1310 -1545 1910
rect -1495 1310 -1445 1910
rect -1395 1310 -1345 1910
rect -1295 1310 -1245 1910
rect -1195 1310 -1145 1910
rect -1095 1310 -1045 1910
rect -995 1310 -945 1910
rect -895 1310 -845 1910
rect -795 1310 -745 1910
rect -695 1310 -645 1910
rect -495 1310 -445 1910
rect -395 1310 -345 1910
rect -295 1310 -245 1910
rect -195 1310 -145 1910
rect -95 1310 -45 1910
rect 5 1310 55 1910
rect 105 1310 155 1910
rect 205 1310 255 1910
rect 305 1310 355 1910
rect 405 1310 455 1910
<< ndiff >>
rect -2345 965 -2295 980
rect -2345 395 -2330 965
rect -2310 395 -2295 965
rect -2345 380 -2295 395
rect -2245 965 -2195 980
rect -2245 395 -2230 965
rect -2210 395 -2195 965
rect -2245 380 -2195 395
rect -2145 965 -2095 980
rect -2145 395 -2130 965
rect -2110 395 -2095 965
rect -2145 380 -2095 395
rect -2045 965 -1995 980
rect -2045 395 -2030 965
rect -2010 395 -1995 965
rect -2045 380 -1995 395
rect -1945 965 -1895 980
rect -1945 395 -1930 965
rect -1910 395 -1895 965
rect -1945 380 -1895 395
rect -1845 965 -1795 980
rect -1845 395 -1830 965
rect -1810 395 -1795 965
rect -1845 380 -1795 395
rect -1745 965 -1695 980
rect -1645 965 -1595 980
rect -1745 395 -1730 965
rect -1710 395 -1695 965
rect -1645 395 -1630 965
rect -1610 395 -1595 965
rect -1745 380 -1695 395
rect -1645 380 -1595 395
rect -1545 965 -1495 980
rect -1545 395 -1530 965
rect -1510 395 -1495 965
rect -1545 380 -1495 395
rect -1445 965 -1395 980
rect -1445 395 -1430 965
rect -1410 395 -1395 965
rect -1445 380 -1395 395
rect -1345 965 -1295 980
rect -1345 395 -1330 965
rect -1310 395 -1295 965
rect -1345 380 -1295 395
rect -1245 965 -1195 980
rect -1245 395 -1230 965
rect -1210 395 -1195 965
rect -1245 380 -1195 395
rect -1145 965 -1095 980
rect -1145 395 -1130 965
rect -1110 395 -1095 965
rect -1145 380 -1095 395
rect -1045 965 -995 980
rect -1045 395 -1030 965
rect -1010 395 -995 965
rect -1045 380 -995 395
rect -945 965 -895 980
rect -945 395 -930 965
rect -910 395 -895 965
rect -945 380 -895 395
rect -845 965 -795 980
rect -845 395 -830 965
rect -810 395 -795 965
rect -845 380 -795 395
rect -745 965 -695 980
rect -745 395 -730 965
rect -710 395 -695 965
rect -745 380 -695 395
rect -645 965 -595 980
rect -545 965 -495 980
rect -645 395 -630 965
rect -610 395 -595 965
rect -545 395 -530 965
rect -510 395 -495 965
rect -645 380 -595 395
rect -545 380 -495 395
rect -445 965 -395 980
rect -445 395 -430 965
rect -410 395 -395 965
rect -445 380 -395 395
rect -345 965 -295 980
rect -345 395 -330 965
rect -310 395 -295 965
rect -345 380 -295 395
rect -245 965 -195 980
rect -245 395 -230 965
rect -210 395 -195 965
rect -245 380 -195 395
rect -145 965 -95 980
rect -145 395 -130 965
rect -110 395 -95 965
rect -145 380 -95 395
rect -45 965 5 980
rect -45 395 -30 965
rect -10 395 5 965
rect -45 380 5 395
rect 55 965 105 980
rect 55 395 70 965
rect 90 395 105 965
rect 55 380 105 395
rect 155 965 205 980
rect 155 395 170 965
rect 190 395 205 965
rect 155 380 205 395
rect 255 965 305 980
rect 255 395 270 965
rect 290 395 305 965
rect 255 380 305 395
rect 355 965 405 980
rect 355 395 370 965
rect 390 395 405 965
rect 355 380 405 395
rect 455 965 505 980
rect 455 395 470 965
rect 490 395 505 965
rect 455 380 505 395
<< pdiff >>
rect -2345 1895 -2295 1910
rect -2345 1325 -2330 1895
rect -2310 1325 -2295 1895
rect -2345 1310 -2295 1325
rect -2245 1895 -2195 1910
rect -2245 1325 -2230 1895
rect -2210 1325 -2195 1895
rect -2245 1310 -2195 1325
rect -2145 1895 -2095 1910
rect -2145 1325 -2130 1895
rect -2110 1325 -2095 1895
rect -2145 1310 -2095 1325
rect -2045 1895 -1995 1910
rect -2045 1325 -2030 1895
rect -2010 1325 -1995 1895
rect -2045 1310 -1995 1325
rect -1945 1895 -1895 1910
rect -1945 1325 -1930 1895
rect -1910 1325 -1895 1895
rect -1945 1310 -1895 1325
rect -1845 1895 -1795 1910
rect -1845 1325 -1830 1895
rect -1810 1325 -1795 1895
rect -1845 1310 -1795 1325
rect -1745 1895 -1695 1910
rect -1645 1895 -1595 1910
rect -1745 1325 -1730 1895
rect -1710 1325 -1695 1895
rect -1645 1325 -1630 1895
rect -1610 1325 -1595 1895
rect -1745 1310 -1695 1325
rect -1645 1310 -1595 1325
rect -1545 1895 -1495 1910
rect -1545 1325 -1530 1895
rect -1510 1325 -1495 1895
rect -1545 1310 -1495 1325
rect -1445 1895 -1395 1910
rect -1445 1325 -1430 1895
rect -1410 1325 -1395 1895
rect -1445 1310 -1395 1325
rect -1345 1895 -1295 1910
rect -1345 1325 -1330 1895
rect -1310 1325 -1295 1895
rect -1345 1310 -1295 1325
rect -1245 1895 -1195 1910
rect -1245 1325 -1230 1895
rect -1210 1325 -1195 1895
rect -1245 1310 -1195 1325
rect -1145 1895 -1095 1910
rect -1145 1325 -1130 1895
rect -1110 1325 -1095 1895
rect -1145 1310 -1095 1325
rect -1045 1895 -995 1910
rect -1045 1325 -1030 1895
rect -1010 1325 -995 1895
rect -1045 1310 -995 1325
rect -945 1895 -895 1910
rect -945 1325 -930 1895
rect -910 1325 -895 1895
rect -945 1310 -895 1325
rect -845 1895 -795 1910
rect -845 1325 -830 1895
rect -810 1325 -795 1895
rect -845 1310 -795 1325
rect -745 1895 -695 1910
rect -745 1325 -730 1895
rect -710 1325 -695 1895
rect -745 1310 -695 1325
rect -645 1895 -595 1910
rect -545 1895 -495 1910
rect -645 1325 -630 1895
rect -610 1325 -595 1895
rect -545 1325 -530 1895
rect -510 1325 -495 1895
rect -645 1310 -595 1325
rect -545 1310 -495 1325
rect -445 1895 -395 1910
rect -445 1325 -430 1895
rect -410 1325 -395 1895
rect -445 1310 -395 1325
rect -345 1895 -295 1910
rect -345 1325 -330 1895
rect -310 1325 -295 1895
rect -345 1310 -295 1325
rect -245 1895 -195 1910
rect -245 1325 -230 1895
rect -210 1325 -195 1895
rect -245 1310 -195 1325
rect -145 1895 -95 1910
rect -145 1325 -130 1895
rect -110 1325 -95 1895
rect -145 1310 -95 1325
rect -45 1895 5 1910
rect -45 1325 -30 1895
rect -10 1325 5 1895
rect -45 1310 5 1325
rect 55 1895 105 1910
rect 55 1325 70 1895
rect 90 1325 105 1895
rect 55 1310 105 1325
rect 155 1895 205 1910
rect 155 1325 170 1895
rect 190 1325 205 1895
rect 155 1310 205 1325
rect 255 1895 305 1910
rect 255 1325 270 1895
rect 290 1325 305 1895
rect 255 1310 305 1325
rect 355 1895 405 1910
rect 355 1325 370 1895
rect 390 1325 405 1895
rect 355 1310 405 1325
rect 455 1895 505 1910
rect 455 1325 470 1895
rect 490 1325 505 1895
rect 455 1310 505 1325
<< ndiffc >>
rect -2330 395 -2310 965
rect -2230 395 -2210 965
rect -2130 395 -2110 965
rect -2030 395 -2010 965
rect -1930 395 -1910 965
rect -1830 395 -1810 965
rect -1730 395 -1710 965
rect -1630 395 -1610 965
rect -1530 395 -1510 965
rect -1430 395 -1410 965
rect -1330 395 -1310 965
rect -1230 395 -1210 965
rect -1130 395 -1110 965
rect -1030 395 -1010 965
rect -930 395 -910 965
rect -830 395 -810 965
rect -730 395 -710 965
rect -630 395 -610 965
rect -530 395 -510 965
rect -430 395 -410 965
rect -330 395 -310 965
rect -230 395 -210 965
rect -130 395 -110 965
rect -30 395 -10 965
rect 70 395 90 965
rect 170 395 190 965
rect 270 395 290 965
rect 370 395 390 965
rect 470 395 490 965
<< pdiffc >>
rect -2330 1325 -2310 1895
rect -2230 1325 -2210 1895
rect -2130 1325 -2110 1895
rect -2030 1325 -2010 1895
rect -1930 1325 -1910 1895
rect -1830 1325 -1810 1895
rect -1730 1325 -1710 1895
rect -1630 1325 -1610 1895
rect -1530 1325 -1510 1895
rect -1430 1325 -1410 1895
rect -1330 1325 -1310 1895
rect -1230 1325 -1210 1895
rect -1130 1325 -1110 1895
rect -1030 1325 -1010 1895
rect -930 1325 -910 1895
rect -830 1325 -810 1895
rect -730 1325 -710 1895
rect -630 1325 -610 1895
rect -530 1325 -510 1895
rect -430 1325 -410 1895
rect -330 1325 -310 1895
rect -230 1325 -210 1895
rect -130 1325 -110 1895
rect -30 1325 -10 1895
rect 70 1325 90 1895
rect 170 1325 190 1895
rect 270 1325 290 1895
rect 370 1325 390 1895
rect 470 1325 490 1895
<< psubdiff >>
rect -2395 965 -2345 980
rect -2395 395 -2380 965
rect -2360 395 -2345 965
rect -2395 380 -2345 395
rect -1695 965 -1645 980
rect -1695 395 -1680 965
rect -1660 395 -1645 965
rect -1695 380 -1645 395
rect -595 965 -545 980
rect -595 395 -580 965
rect -560 395 -545 965
rect -595 380 -545 395
rect 505 965 555 980
rect 505 395 520 965
rect 540 395 555 965
rect 505 380 555 395
<< nsubdiff >>
rect -2395 1895 -2345 1910
rect -2395 1325 -2380 1895
rect -2360 1325 -2345 1895
rect -2395 1310 -2345 1325
rect -1695 1895 -1645 1910
rect -1695 1325 -1680 1895
rect -1660 1325 -1645 1895
rect -1695 1310 -1645 1325
rect -595 1895 -545 1910
rect -595 1325 -580 1895
rect -560 1325 -545 1895
rect -595 1310 -545 1325
rect 505 1895 555 1910
rect 505 1325 520 1895
rect 540 1325 555 1895
rect 505 1310 555 1325
<< psubdiffcont >>
rect -2380 395 -2360 965
rect -1680 395 -1660 965
rect -580 395 -560 965
rect 520 395 540 965
<< nsubdiffcont >>
rect -2380 1325 -2360 1895
rect -1680 1325 -1660 1895
rect -580 1325 -560 1895
rect 520 1325 540 1895
<< poly >>
rect -2295 1955 -2245 1970
rect -2295 1935 -2280 1955
rect -2260 1935 -2245 1955
rect -2295 1910 -2245 1935
rect -1795 1955 -1745 1970
rect -1795 1935 -1780 1955
rect -1760 1935 -1745 1955
rect -2195 1910 -2145 1925
rect -2095 1910 -2045 1925
rect -1995 1910 -1945 1925
rect -1895 1910 -1845 1925
rect -1795 1910 -1745 1935
rect -1495 1955 -745 2005
rect -1595 1910 -1545 1925
rect -1495 1910 -1445 1955
rect -1395 1910 -1345 1955
rect -1295 1910 -1245 1955
rect -1195 1910 -1145 1925
rect -1095 1910 -1045 1925
rect -995 1910 -945 1955
rect -895 1910 -845 1955
rect -795 1910 -745 1955
rect -495 1955 -445 1970
rect -495 1935 -480 1955
rect -460 1935 -445 1955
rect -695 1910 -645 1925
rect -495 1910 -445 1935
rect 405 1955 455 1970
rect 405 1935 420 1955
rect 440 1935 455 1955
rect -395 1910 -345 1925
rect -295 1910 -245 1925
rect -195 1910 -145 1925
rect -95 1910 -45 1925
rect 5 1910 55 1925
rect 105 1910 155 1925
rect 205 1910 255 1925
rect 305 1910 355 1925
rect 405 1910 455 1935
rect -2295 1295 -2245 1310
rect -2195 1275 -2145 1310
rect -2195 1255 -2180 1275
rect -2160 1255 -2145 1275
rect -2195 1240 -2145 1255
rect -2095 1295 -2045 1310
rect -1995 1295 -1945 1310
rect -2095 1280 -1945 1295
rect -2095 1260 -2030 1280
rect -2010 1260 -1945 1280
rect -2095 1245 -1945 1260
rect -1895 1275 -1845 1310
rect -1795 1295 -1745 1310
rect -1895 1255 -1880 1275
rect -1860 1255 -1845 1275
rect -1895 1240 -1845 1255
rect -1595 1285 -1545 1310
rect -1595 1265 -1580 1285
rect -1560 1265 -1545 1285
rect -1595 1250 -1545 1265
rect -1495 1295 -1445 1310
rect -1395 1295 -1345 1310
rect -1295 1295 -1245 1310
rect -1495 1285 -1245 1295
rect -1495 1265 -1380 1285
rect -1360 1265 -1245 1285
rect -1495 1245 -1245 1265
rect -1195 1295 -1145 1310
rect -1095 1295 -1045 1310
rect -1195 1285 -1045 1295
rect -1195 1265 -1130 1285
rect -1110 1265 -1045 1285
rect -1195 1245 -1045 1265
rect -995 1295 -945 1310
rect -895 1295 -845 1310
rect -795 1295 -745 1310
rect -995 1285 -745 1295
rect -995 1265 -880 1285
rect -860 1265 -745 1285
rect -995 1235 -745 1265
rect -695 1285 -645 1310
rect -495 1295 -445 1310
rect -395 1295 -345 1310
rect -295 1295 -245 1310
rect -195 1295 -145 1310
rect -95 1295 -45 1310
rect 5 1295 55 1310
rect 105 1295 155 1310
rect 205 1295 255 1310
rect 305 1295 355 1310
rect 405 1295 455 1310
rect -695 1265 -680 1285
rect -660 1265 -645 1285
rect -695 1250 -645 1265
rect -395 1275 355 1295
rect -395 1255 -230 1275
rect -210 1255 170 1275
rect 190 1255 355 1275
rect -395 1245 355 1255
rect -2195 1035 -1845 1045
rect -2195 1015 -2130 1035
rect -2110 1015 -1930 1035
rect -1910 1015 -1845 1035
rect -2195 995 -1845 1015
rect -1495 1035 -745 1045
rect -1495 1015 -1330 1035
rect -1310 1015 -930 1035
rect -910 1015 -745 1035
rect -1495 995 -745 1015
rect -495 1025 -445 1040
rect -495 1005 -480 1025
rect -460 1005 -445 1025
rect -2295 980 -2245 995
rect -2195 980 -2145 995
rect -2095 980 -2045 995
rect -1995 980 -1945 995
rect -1895 980 -1845 995
rect -1795 980 -1745 995
rect -1595 980 -1545 995
rect -1495 980 -1445 995
rect -1395 980 -1345 995
rect -1295 980 -1245 995
rect -1195 980 -1145 995
rect -1095 980 -1045 995
rect -995 980 -945 995
rect -895 980 -845 995
rect -795 980 -745 995
rect -695 980 -645 995
rect -495 980 -445 1005
rect -395 1035 -145 1045
rect -395 1015 -280 1035
rect -260 1015 -145 1035
rect -395 995 -145 1015
rect -395 980 -345 995
rect -295 980 -245 995
rect -195 980 -145 995
rect -95 1035 55 1045
rect -95 1015 -30 1035
rect -10 1015 55 1035
rect -95 1000 55 1015
rect -95 980 -45 1000
rect 5 980 55 1000
rect 105 1035 355 1045
rect 105 1015 220 1035
rect 240 1015 355 1035
rect 105 1005 355 1015
rect 105 980 155 1005
rect 205 980 255 1005
rect 305 980 355 1005
rect 405 1030 455 1045
rect 405 1010 420 1030
rect 440 1010 455 1030
rect 405 980 455 1010
rect -2295 355 -2245 380
rect -2195 365 -2145 380
rect -2095 365 -2045 380
rect -1995 365 -1945 380
rect -1895 365 -1845 380
rect -2295 335 -2280 355
rect -2260 335 -2245 355
rect -2295 320 -2245 335
rect -1795 355 -1745 380
rect -1795 335 -1780 355
rect -1760 335 -1745 355
rect -1795 320 -1745 335
rect -1595 355 -1545 380
rect -1495 365 -1445 380
rect -1395 365 -1345 380
rect -1295 365 -1245 380
rect -1195 365 -1145 380
rect -1095 365 -1045 380
rect -995 365 -945 380
rect -895 365 -845 380
rect -795 365 -745 380
rect -1595 335 -1580 355
rect -1560 335 -1545 355
rect -1595 320 -1545 335
rect -695 355 -645 380
rect -495 365 -445 380
rect -695 335 -680 355
rect -660 335 -645 355
rect -695 320 -645 335
rect -395 335 -345 380
rect -295 335 -245 380
rect -195 335 -145 380
rect -95 365 -45 380
rect 5 365 55 380
rect 105 335 155 380
rect 205 335 255 380
rect 305 335 355 380
rect 405 365 455 380
rect -395 285 355 335
<< polycont >>
rect -2280 1935 -2260 1955
rect -1780 1935 -1760 1955
rect -480 1935 -460 1955
rect 420 1935 440 1955
rect -2180 1255 -2160 1275
rect -2030 1260 -2010 1280
rect -1880 1255 -1860 1275
rect -1580 1265 -1560 1285
rect -1380 1265 -1360 1285
rect -1130 1265 -1110 1285
rect -880 1265 -860 1285
rect -680 1265 -660 1285
rect -230 1255 -210 1275
rect 170 1255 190 1275
rect -2130 1015 -2110 1035
rect -1930 1015 -1910 1035
rect -1330 1015 -1310 1035
rect -930 1015 -910 1035
rect -480 1005 -460 1025
rect -280 1015 -260 1035
rect -30 1015 -10 1035
rect 220 1015 240 1035
rect 420 1010 440 1030
rect -2280 335 -2260 355
rect -1780 335 -1760 355
rect -1580 335 -1560 355
rect -680 335 -660 355
<< locali >>
rect -2390 1955 -2250 1965
rect -2390 1935 -2280 1955
rect -2260 1935 -2250 1955
rect -2390 1925 -2250 1935
rect -1790 1955 -1650 1965
rect -1790 1935 -1780 1955
rect -1760 1935 -1650 1955
rect -1790 1925 -1650 1935
rect -2390 1895 -2300 1925
rect -1740 1905 -1650 1925
rect -1440 1925 -800 1965
rect -2390 1325 -2380 1895
rect -2360 1325 -2330 1895
rect -2310 1325 -2300 1895
rect -2390 1315 -2300 1325
rect -2240 1895 -2200 1905
rect -2240 1325 -2230 1895
rect -2210 1325 -2200 1895
rect -2240 1285 -2200 1325
rect -2140 1895 -2100 1905
rect -2140 1325 -2130 1895
rect -2110 1325 -2100 1895
rect -2140 1315 -2100 1325
rect -2040 1895 -2000 1905
rect -2040 1325 -2030 1895
rect -2010 1325 -2000 1895
rect -2040 1295 -2000 1325
rect -1940 1895 -1900 1905
rect -1940 1325 -1930 1895
rect -1910 1325 -1900 1895
rect -1940 1315 -1900 1325
rect -1840 1895 -1800 1905
rect -1840 1325 -1830 1895
rect -1810 1325 -1800 1895
rect -2240 1275 -2150 1285
rect -2240 1255 -2180 1275
rect -2160 1255 -2150 1275
rect -2240 1245 -2150 1255
rect -2045 1280 -1995 1295
rect -1840 1285 -1800 1325
rect -1740 1895 -1600 1905
rect -1740 1325 -1730 1895
rect -1710 1325 -1680 1895
rect -1660 1325 -1630 1895
rect -1610 1325 -1600 1895
rect -1740 1315 -1600 1325
rect -1540 1895 -1500 1905
rect -1540 1325 -1530 1895
rect -1510 1325 -1500 1895
rect -1540 1315 -1500 1325
rect -1440 1895 -1400 1925
rect -1440 1325 -1430 1895
rect -1410 1325 -1400 1895
rect -1440 1315 -1400 1325
rect -1340 1895 -1300 1905
rect -1340 1325 -1330 1895
rect -1310 1325 -1300 1895
rect -1340 1315 -1300 1325
rect -1240 1895 -1200 1925
rect -1240 1325 -1230 1895
rect -1210 1325 -1200 1895
rect -1240 1315 -1200 1325
rect -1140 1895 -1100 1905
rect -1140 1325 -1130 1895
rect -1110 1325 -1100 1895
rect -2045 1260 -2030 1280
rect -2010 1260 -1995 1280
rect -2045 1245 -1995 1260
rect -1890 1275 -1800 1285
rect -1890 1255 -1880 1275
rect -1860 1255 -1800 1275
rect -1690 1295 -1600 1315
rect -1690 1285 -1550 1295
rect -1690 1265 -1580 1285
rect -1560 1265 -1550 1285
rect -1690 1255 -1550 1265
rect -1390 1285 -1350 1295
rect -1390 1265 -1380 1285
rect -1360 1265 -1350 1285
rect -1890 1245 -1800 1255
rect -2390 965 -2300 975
rect -2390 395 -2380 965
rect -2360 395 -2330 965
rect -2310 395 -2300 965
rect -2390 365 -2300 395
rect -2240 965 -2200 1245
rect -2140 1035 -1900 1045
rect -2140 1015 -2130 1035
rect -2110 1015 -1930 1035
rect -1910 1015 -1900 1035
rect -2140 1005 -1900 1015
rect -2240 395 -2230 965
rect -2210 395 -2200 965
rect -2240 385 -2200 395
rect -2140 965 -2100 975
rect -2140 395 -2130 965
rect -2110 395 -2100 965
rect -2140 385 -2100 395
rect -2040 965 -2000 1005
rect -2040 395 -2030 965
rect -2010 395 -2000 965
rect -2040 385 -2000 395
rect -1940 965 -1900 975
rect -1940 395 -1930 965
rect -1910 395 -1900 965
rect -1940 385 -1900 395
rect -1840 965 -1800 1245
rect -1390 1190 -1350 1265
rect -1540 1150 -1350 1190
rect -1140 1285 -1100 1325
rect -1040 1895 -1000 1925
rect -1040 1325 -1030 1895
rect -1010 1325 -1000 1895
rect -1040 1315 -1000 1325
rect -940 1895 -900 1905
rect -940 1325 -930 1895
rect -910 1325 -900 1895
rect -940 1315 -900 1325
rect -840 1895 -800 1925
rect -590 1955 -450 1965
rect -590 1935 -480 1955
rect -460 1935 -450 1955
rect -590 1925 -450 1935
rect 410 1955 550 1965
rect 410 1935 420 1955
rect 440 1935 550 1955
rect 410 1925 550 1935
rect -590 1905 -500 1925
rect -840 1325 -830 1895
rect -810 1325 -800 1895
rect -840 1315 -800 1325
rect -740 1895 -700 1905
rect -740 1325 -730 1895
rect -710 1325 -700 1895
rect -740 1315 -700 1325
rect -640 1895 -500 1905
rect -640 1325 -630 1895
rect -610 1325 -580 1895
rect -560 1325 -530 1895
rect -510 1325 -500 1895
rect -640 1315 -500 1325
rect -440 1895 -400 1905
rect -440 1325 -430 1895
rect -410 1325 -400 1895
rect -640 1295 -550 1315
rect -1140 1265 -1130 1285
rect -1110 1265 -1100 1285
rect -1140 1210 -1100 1265
rect -890 1285 -850 1295
rect -890 1265 -880 1285
rect -860 1265 -850 1285
rect -1140 1200 -1090 1210
rect -1140 1170 -1130 1200
rect -1100 1170 -1090 1200
rect -1140 1160 -1090 1170
rect -890 1190 -850 1265
rect -690 1285 -550 1295
rect -690 1265 -680 1285
rect -660 1265 -550 1285
rect -690 1255 -550 1265
rect -440 1195 -400 1325
rect -340 1895 -300 1905
rect -340 1325 -330 1895
rect -310 1325 -300 1895
rect -340 1315 -300 1325
rect -240 1895 -200 1905
rect -240 1325 -230 1895
rect -210 1325 -200 1895
rect -240 1315 -200 1325
rect -140 1895 -100 1905
rect -140 1325 -130 1895
rect -110 1325 -100 1895
rect -140 1315 -100 1325
rect -40 1895 0 1905
rect -40 1325 -30 1895
rect -10 1325 0 1895
rect -240 1275 -200 1285
rect -240 1255 -230 1275
rect -210 1255 -200 1275
rect -240 1245 -200 1255
rect -1840 395 -1830 965
rect -1810 395 -1800 965
rect -1840 385 -1800 395
rect -1740 965 -1600 975
rect -1740 395 -1730 965
rect -1710 395 -1680 965
rect -1660 395 -1630 965
rect -1610 395 -1600 965
rect -1740 365 -1600 395
rect -1540 965 -1500 1150
rect -1340 1035 -1300 1045
rect -1340 1015 -1330 1035
rect -1310 1015 -1300 1035
rect -1340 1005 -1300 1015
rect -1540 395 -1530 965
rect -1510 395 -1500 965
rect -1540 385 -1500 395
rect -1440 965 -1400 975
rect -1440 395 -1430 965
rect -1410 395 -1400 965
rect -1440 385 -1400 395
rect -1340 965 -1300 975
rect -1340 395 -1330 965
rect -1310 395 -1300 965
rect -1340 385 -1300 395
rect -1240 965 -1200 975
rect -1240 395 -1230 965
rect -1210 395 -1200 965
rect -1240 385 -1200 395
rect -1140 965 -1100 1160
rect -890 1150 -700 1190
rect -440 1155 -250 1195
rect -940 1035 -900 1045
rect -940 1015 -930 1035
rect -910 1015 -900 1035
rect -940 1005 -900 1015
rect -1140 395 -1130 965
rect -1110 395 -1100 965
rect -1140 385 -1100 395
rect -1040 965 -1000 975
rect -1040 395 -1030 965
rect -1010 395 -1000 965
rect -1040 385 -1000 395
rect -940 965 -900 975
rect -940 395 -930 965
rect -910 395 -900 965
rect -940 385 -900 395
rect -840 965 -800 975
rect -840 395 -830 965
rect -810 395 -800 965
rect -840 385 -800 395
rect -740 965 -700 1150
rect -290 1035 -250 1155
rect -590 1025 -450 1035
rect -590 1005 -480 1025
rect -460 1005 -450 1025
rect -290 1015 -280 1035
rect -260 1015 -250 1035
rect -290 1005 -250 1015
rect -40 1135 0 1325
rect 60 1895 100 1905
rect 60 1325 70 1895
rect 90 1325 100 1895
rect 60 1315 100 1325
rect 160 1895 200 1905
rect 160 1325 170 1895
rect 190 1325 200 1895
rect 160 1315 200 1325
rect 260 1895 300 1905
rect 260 1325 270 1895
rect 290 1325 300 1895
rect 260 1315 300 1325
rect 360 1895 400 1905
rect 360 1325 370 1895
rect 390 1325 400 1895
rect 160 1275 200 1285
rect 160 1255 170 1275
rect 190 1255 200 1275
rect 160 1245 200 1255
rect 360 1195 400 1325
rect 460 1895 550 1925
rect 460 1325 470 1895
rect 490 1325 520 1895
rect 540 1325 550 1895
rect 460 1315 550 1325
rect 210 1155 400 1195
rect -40 1125 10 1135
rect -40 1095 -30 1125
rect 0 1095 10 1125
rect -40 1085 10 1095
rect -40 1035 0 1085
rect -40 1015 -30 1035
rect -10 1015 0 1035
rect -590 995 -450 1005
rect -590 975 -500 995
rect -740 395 -730 965
rect -710 395 -700 965
rect -740 385 -700 395
rect -640 965 -500 975
rect -640 395 -630 965
rect -610 395 -580 965
rect -560 395 -530 965
rect -510 395 -500 965
rect -640 385 -500 395
rect -440 965 -400 975
rect -440 395 -430 965
rect -410 395 -400 965
rect -440 385 -400 395
rect -340 965 -300 975
rect -340 395 -330 965
rect -310 395 -300 965
rect -640 365 -550 385
rect -2390 355 -2250 365
rect -2390 335 -2280 355
rect -2260 335 -2250 355
rect -2390 325 -2250 335
rect -1790 355 -1550 365
rect -1790 335 -1780 355
rect -1760 335 -1580 355
rect -1560 335 -1550 355
rect -1790 325 -1550 335
rect -690 355 -550 365
rect -690 335 -680 355
rect -660 335 -550 355
rect -690 325 -550 335
rect -340 365 -300 395
rect -240 965 -200 975
rect -240 395 -230 965
rect -210 395 -200 965
rect -240 385 -200 395
rect -140 965 -100 975
rect -140 395 -130 965
rect -110 395 -100 965
rect -140 365 -100 395
rect -40 965 0 1015
rect 210 1035 250 1155
rect 210 1015 220 1035
rect 240 1015 250 1035
rect 210 1005 250 1015
rect 410 1030 550 1040
rect 410 1010 420 1030
rect 440 1010 550 1030
rect 410 1000 550 1010
rect -40 395 -30 965
rect -10 395 0 965
rect -40 385 0 395
rect 60 965 100 975
rect 60 395 70 965
rect 90 395 100 965
rect 60 365 100 395
rect 160 965 200 975
rect 160 395 170 965
rect 190 395 200 965
rect 160 385 200 395
rect 260 965 300 975
rect 260 395 270 965
rect 290 395 300 965
rect 260 365 300 395
rect 360 965 400 975
rect 360 395 370 965
rect 390 395 400 965
rect 360 385 400 395
rect 460 965 550 1000
rect 460 395 470 965
rect 490 395 520 965
rect 540 395 550 965
rect 460 385 550 395
rect -340 325 300 365
<< viali >>
rect -2380 1325 -2360 1895
rect -2330 1325 -2310 1895
rect -2130 1325 -2110 1895
rect -2030 1325 -2010 1895
rect -1930 1325 -1910 1895
rect -2180 1255 -2160 1275
rect -1730 1325 -1710 1895
rect -1680 1325 -1660 1895
rect -1630 1325 -1610 1895
rect -1530 1325 -1510 1895
rect -1880 1255 -1860 1275
rect -2380 395 -2360 965
rect -2330 395 -2310 965
rect -2130 1015 -2110 1035
rect -1930 1015 -1910 1035
rect -2130 395 -2110 965
rect -1930 395 -1910 965
rect -730 1325 -710 1895
rect -630 1325 -610 1895
rect -580 1325 -560 1895
rect -530 1325 -510 1895
rect -1130 1170 -1100 1200
rect -130 1325 -110 1895
rect -230 1255 -210 1275
rect -1730 395 -1710 965
rect -1680 395 -1660 965
rect -1630 395 -1610 965
rect -1330 1015 -1310 1035
rect -1230 395 -1210 965
rect -930 1015 -910 1035
rect -1030 395 -1010 965
rect 70 1325 90 1895
rect 170 1255 190 1275
rect 470 1325 490 1895
rect 520 1325 540 1895
rect -30 1095 0 1125
rect -630 395 -610 965
rect -580 395 -560 965
rect -530 395 -510 965
rect -430 395 -410 965
rect 370 395 390 965
rect 470 395 490 965
rect 520 395 540 965
<< metal1 >>
rect -2395 1895 560 1905
rect -2395 1325 -2380 1895
rect -2360 1325 -2330 1895
rect -2310 1325 -2130 1895
rect -2110 1325 -2030 1895
rect -2010 1325 -1930 1895
rect -1910 1325 -1730 1895
rect -1710 1325 -1680 1895
rect -1660 1325 -1630 1895
rect -1610 1325 -1530 1895
rect -1510 1325 -730 1895
rect -710 1325 -630 1895
rect -610 1325 -580 1895
rect -560 1325 -530 1895
rect -510 1325 -130 1895
rect -110 1325 70 1895
rect 90 1325 470 1895
rect 490 1325 520 1895
rect 540 1325 560 1895
rect -2395 1315 560 1325
rect -2195 1275 555 1285
rect -2195 1255 -2180 1275
rect -2160 1255 -1880 1275
rect -1860 1255 -230 1275
rect -210 1255 170 1275
rect 190 1255 555 1275
rect -2195 1235 555 1255
rect -1140 1200 555 1210
rect -1140 1170 -1130 1200
rect -1100 1170 555 1200
rect -2400 1115 -1995 1165
rect -1140 1160 555 1170
rect -2045 1055 -1995 1115
rect -40 1125 555 1135
rect -40 1095 -30 1125
rect 0 1095 555 1125
rect -40 1085 555 1095
rect -2195 1035 555 1055
rect -2195 1015 -2130 1035
rect -2110 1015 -1930 1035
rect -1910 1015 -1330 1035
rect -1310 1015 -930 1035
rect -910 1015 555 1035
rect -2195 1005 555 1015
rect -2400 965 555 975
rect -2400 395 -2380 965
rect -2360 395 -2330 965
rect -2310 395 -2130 965
rect -2110 395 -1930 965
rect -1910 395 -1730 965
rect -1710 395 -1680 965
rect -1660 395 -1630 965
rect -1610 395 -1230 965
rect -1210 395 -1030 965
rect -1010 395 -630 965
rect -610 395 -580 965
rect -560 395 -530 965
rect -510 395 -430 965
rect -410 395 370 965
rect 390 395 470 965
rect 490 395 520 965
rect 540 395 555 965
rect -2400 385 555 395
<< labels >>
rlabel metal1 555 1260 555 1260 3 Vbp
rlabel metal1 555 1185 555 1185 3 Vcp
rlabel metal1 555 1110 555 1110 3 Vcn
rlabel metal1 555 1030 555 1030 3 Vbn
rlabel metal1 -2400 680 -2400 680 7 GND
rlabel metal1 -2395 1610 -2395 1610 7 VDD
rlabel ndiff -1325 980 -1325 980 1 net2
<< end >>
