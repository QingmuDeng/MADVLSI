magic
tech sky130A
timestamp 1615258659
<< nmos >>
rect -2295 315 -2245 915
rect -2195 315 -2145 915
rect -2095 315 -2045 915
rect -1995 315 -1945 915
rect -1895 315 -1845 915
rect -1795 315 -1745 915
rect -1595 315 -1545 915
rect -1495 315 -1445 915
rect -1395 315 -1345 915
rect -1295 315 -1245 915
rect -1195 315 -1145 915
rect -1095 315 -1045 915
rect -995 315 -945 915
rect -895 315 -845 915
rect -795 315 -745 915
rect -695 315 -645 915
rect -495 315 -445 915
rect -395 315 -345 915
rect -295 315 -245 915
rect -195 315 -145 915
rect -95 315 -45 915
rect 5 315 55 915
rect 105 315 155 915
rect 205 315 255 915
rect 305 315 355 915
rect 405 315 455 915
<< ndiff >>
rect -2345 900 -2295 915
rect -2345 330 -2330 900
rect -2310 330 -2295 900
rect -2345 315 -2295 330
rect -2245 900 -2195 915
rect -2245 330 -2230 900
rect -2210 330 -2195 900
rect -2245 315 -2195 330
rect -2145 900 -2095 915
rect -2145 330 -2130 900
rect -2110 330 -2095 900
rect -2145 315 -2095 330
rect -2045 900 -1995 915
rect -2045 330 -2030 900
rect -2010 330 -1995 900
rect -2045 315 -1995 330
rect -1945 900 -1895 915
rect -1945 330 -1930 900
rect -1910 330 -1895 900
rect -1945 315 -1895 330
rect -1845 900 -1795 915
rect -1845 330 -1830 900
rect -1810 330 -1795 900
rect -1845 315 -1795 330
rect -1745 900 -1695 915
rect -1645 900 -1595 915
rect -1745 330 -1730 900
rect -1710 330 -1695 900
rect -1645 330 -1630 900
rect -1610 330 -1595 900
rect -1745 315 -1695 330
rect -1645 315 -1595 330
rect -1545 900 -1495 915
rect -1545 330 -1530 900
rect -1510 330 -1495 900
rect -1545 315 -1495 330
rect -1445 900 -1395 915
rect -1445 330 -1430 900
rect -1410 330 -1395 900
rect -1445 315 -1395 330
rect -1345 900 -1295 915
rect -1345 330 -1330 900
rect -1310 330 -1295 900
rect -1345 315 -1295 330
rect -1245 900 -1195 915
rect -1245 330 -1230 900
rect -1210 330 -1195 900
rect -1245 315 -1195 330
rect -1145 900 -1095 915
rect -1145 330 -1130 900
rect -1110 330 -1095 900
rect -1145 315 -1095 330
rect -1045 900 -995 915
rect -1045 330 -1030 900
rect -1010 330 -995 900
rect -1045 315 -995 330
rect -945 900 -895 915
rect -945 330 -930 900
rect -910 330 -895 900
rect -945 315 -895 330
rect -845 900 -795 915
rect -845 330 -830 900
rect -810 330 -795 900
rect -845 315 -795 330
rect -745 900 -695 915
rect -745 330 -730 900
rect -710 330 -695 900
rect -745 315 -695 330
rect -645 900 -595 915
rect -545 900 -495 915
rect -645 330 -630 900
rect -610 330 -595 900
rect -545 330 -530 900
rect -510 330 -495 900
rect -645 315 -595 330
rect -545 315 -495 330
rect -445 900 -395 915
rect -445 330 -430 900
rect -410 330 -395 900
rect -445 315 -395 330
rect -345 900 -295 915
rect -345 330 -330 900
rect -310 330 -295 900
rect -345 315 -295 330
rect -245 900 -195 915
rect -245 330 -230 900
rect -210 330 -195 900
rect -245 315 -195 330
rect -145 900 -95 915
rect -145 330 -130 900
rect -110 330 -95 900
rect -145 315 -95 330
rect -45 900 5 915
rect -45 330 -30 900
rect -10 330 5 900
rect -45 315 5 330
rect 55 900 105 915
rect 55 330 70 900
rect 90 330 105 900
rect 55 315 105 330
rect 155 900 205 915
rect 155 330 170 900
rect 190 330 205 900
rect 155 315 205 330
rect 255 900 305 915
rect 255 330 270 900
rect 290 330 305 900
rect 255 315 305 330
rect 355 900 405 915
rect 355 330 370 900
rect 390 330 405 900
rect 355 315 405 330
rect 455 900 505 915
rect 455 330 470 900
rect 490 330 505 900
rect 455 315 505 330
<< ndiffc >>
rect -2330 330 -2310 900
rect -2230 330 -2210 900
rect -2130 330 -2110 900
rect -2030 330 -2010 900
rect -1930 330 -1910 900
rect -1830 330 -1810 900
rect -1730 330 -1710 900
rect -1630 330 -1610 900
rect -1530 330 -1510 900
rect -1430 330 -1410 900
rect -1330 330 -1310 900
rect -1230 330 -1210 900
rect -1130 330 -1110 900
rect -1030 330 -1010 900
rect -930 330 -910 900
rect -830 330 -810 900
rect -730 330 -710 900
rect -630 330 -610 900
rect -530 330 -510 900
rect -430 330 -410 900
rect -330 330 -310 900
rect -230 330 -210 900
rect -130 330 -110 900
rect -30 330 -10 900
rect 70 330 90 900
rect 170 330 190 900
rect 270 330 290 900
rect 370 330 390 900
rect 470 330 490 900
<< psubdiff >>
rect -2395 900 -2345 915
rect -2395 330 -2380 900
rect -2360 330 -2345 900
rect -2395 315 -2345 330
rect -1695 900 -1645 915
rect -1695 330 -1680 900
rect -1660 330 -1645 900
rect -1695 315 -1645 330
rect -595 900 -545 915
rect -595 330 -580 900
rect -560 330 -545 900
rect -595 315 -545 330
rect 505 900 555 915
rect 505 330 520 900
rect 540 330 555 900
rect 505 315 555 330
<< psubdiffcont >>
rect -2380 330 -2360 900
rect -1680 330 -1660 900
rect -580 330 -560 900
rect 520 330 540 900
<< poly >>
rect -2295 915 -2245 930
rect -2195 915 -2145 930
rect -2095 915 -2045 930
rect -1995 915 -1945 930
rect -1895 915 -1845 930
rect -1795 915 -1745 930
rect -1595 915 -1545 930
rect -1495 915 -1445 930
rect -1395 915 -1345 930
rect -1295 915 -1245 930
rect -1195 915 -1145 930
rect -1095 915 -1045 930
rect -995 915 -945 930
rect -895 915 -845 930
rect -795 915 -745 930
rect -695 915 -645 930
rect -495 915 -445 930
rect -395 915 -345 930
rect -295 915 -245 930
rect -195 915 -145 930
rect -95 915 -45 930
rect 5 915 55 930
rect 105 915 155 930
rect 205 915 255 930
rect 305 915 355 930
rect 405 915 455 930
rect -2295 300 -2245 315
rect -2195 300 -2145 315
rect -2095 300 -2045 315
rect -1995 300 -1945 315
rect -1895 300 -1845 315
rect -1795 300 -1745 315
rect -1595 300 -1545 315
rect -1495 300 -1445 315
rect -1395 300 -1345 315
rect -1295 300 -1245 315
rect -1195 300 -1145 315
rect -1095 300 -1045 315
rect -995 300 -945 315
rect -895 300 -845 315
rect -795 300 -745 315
rect -695 300 -645 315
rect -495 300 -445 315
rect -395 300 -345 315
rect -295 300 -245 315
rect -195 300 -145 315
rect -95 300 -45 315
rect 5 300 55 315
rect 105 300 155 315
rect 205 300 255 315
rect 305 300 355 315
rect 405 300 455 315
<< locali >>
rect -2390 900 -2300 910
rect -2390 330 -2380 900
rect -2360 330 -2330 900
rect -2310 330 -2300 900
rect -2390 320 -2300 330
rect -2240 900 -2200 910
rect -2240 330 -2230 900
rect -2210 330 -2200 900
rect -2240 320 -2200 330
rect -2140 900 -2100 910
rect -2140 330 -2130 900
rect -2110 330 -2100 900
rect -2140 320 -2100 330
rect -2040 900 -2000 910
rect -2040 330 -2030 900
rect -2010 330 -2000 900
rect -2040 320 -2000 330
rect -1940 900 -1900 910
rect -1940 330 -1930 900
rect -1910 330 -1900 900
rect -1940 320 -1900 330
rect -1840 900 -1800 910
rect -1840 330 -1830 900
rect -1810 330 -1800 900
rect -1840 320 -1800 330
rect -1740 900 -1600 910
rect -1740 330 -1730 900
rect -1710 330 -1680 900
rect -1660 330 -1630 900
rect -1610 330 -1600 900
rect -1740 320 -1600 330
rect -1540 900 -1500 910
rect -1540 330 -1530 900
rect -1510 330 -1500 900
rect -1540 320 -1500 330
rect -1440 900 -1400 910
rect -1440 330 -1430 900
rect -1410 330 -1400 900
rect -1440 320 -1400 330
rect -1340 900 -1300 910
rect -1340 330 -1330 900
rect -1310 330 -1300 900
rect -1340 320 -1300 330
rect -1240 900 -1200 910
rect -1240 330 -1230 900
rect -1210 330 -1200 900
rect -1240 320 -1200 330
rect -1140 900 -1100 910
rect -1140 330 -1130 900
rect -1110 330 -1100 900
rect -1140 320 -1100 330
rect -1040 900 -1000 910
rect -1040 330 -1030 900
rect -1010 330 -1000 900
rect -1040 320 -1000 330
rect -940 900 -900 910
rect -940 330 -930 900
rect -910 330 -900 900
rect -940 320 -900 330
rect -840 900 -800 910
rect -840 330 -830 900
rect -810 330 -800 900
rect -840 320 -800 330
rect -740 900 -700 910
rect -740 330 -730 900
rect -710 330 -700 900
rect -740 320 -700 330
rect -640 900 -500 910
rect -640 330 -630 900
rect -610 330 -580 900
rect -560 330 -530 900
rect -510 330 -500 900
rect -640 320 -500 330
rect -440 900 -400 910
rect -440 330 -430 900
rect -410 330 -400 900
rect -440 320 -400 330
rect -340 900 -300 910
rect -340 330 -330 900
rect -310 330 -300 900
rect -340 320 -300 330
rect -240 900 -200 910
rect -240 330 -230 900
rect -210 330 -200 900
rect -240 320 -200 330
rect -140 900 -100 910
rect -140 330 -130 900
rect -110 330 -100 900
rect -140 320 -100 330
rect -40 900 0 910
rect -40 330 -30 900
rect -10 330 0 900
rect -40 320 0 330
rect 60 900 100 910
rect 60 330 70 900
rect 90 330 100 900
rect 60 320 100 330
rect 160 900 200 910
rect 160 330 170 900
rect 190 330 200 900
rect 160 320 200 330
rect 260 900 300 910
rect 260 330 270 900
rect 290 330 300 900
rect 260 320 300 330
rect 360 900 400 910
rect 360 330 370 900
rect 390 330 400 900
rect 360 320 400 330
rect 460 900 550 910
rect 460 330 470 900
rect 490 330 520 900
rect 540 330 550 900
rect 460 320 550 330
<< end >>
