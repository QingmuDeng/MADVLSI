magic
tech sky130A
timestamp 1614043687
<< nwell >>
rect -85 195 255 610
<< nmos >>
rect 0 60 15 160
rect 40 60 55 160
rect 105 60 120 160
rect 170 60 185 160
rect 0 -215 15 -115
rect 40 -215 55 -115
rect 105 -215 120 -115
rect 170 -215 185 -115
<< pmos >>
rect 0 490 15 590
rect 65 490 80 590
rect 130 490 145 590
rect 170 490 185 590
rect 0 215 15 315
rect 65 215 80 315
rect 130 215 145 315
rect 170 215 185 315
<< ndiff >>
rect -50 145 0 160
rect -50 75 -35 145
rect -15 75 0 145
rect -50 60 0 75
rect 15 60 40 160
rect 55 145 105 160
rect 55 75 70 145
rect 90 75 105 145
rect 55 60 105 75
rect 120 145 170 160
rect 120 75 135 145
rect 155 75 170 145
rect 120 60 170 75
rect 185 145 235 160
rect 185 75 200 145
rect 220 75 235 145
rect 185 60 235 75
rect -50 -130 0 -115
rect -50 -200 -35 -130
rect -15 -200 0 -130
rect -50 -215 0 -200
rect 15 -215 40 -115
rect 55 -130 105 -115
rect 55 -200 70 -130
rect 90 -200 105 -130
rect 55 -215 105 -200
rect 120 -130 170 -115
rect 120 -200 135 -130
rect 155 -200 170 -130
rect 120 -215 170 -200
rect 185 -130 235 -115
rect 185 -200 200 -130
rect 220 -200 235 -130
rect 185 -215 235 -200
<< pdiff >>
rect -50 575 0 590
rect -50 505 -35 575
rect -15 505 0 575
rect -50 490 0 505
rect 15 575 65 590
rect 15 505 30 575
rect 50 505 65 575
rect 15 490 65 505
rect 80 575 130 590
rect 80 505 95 575
rect 115 505 130 575
rect 80 490 130 505
rect 145 490 170 590
rect 185 575 235 590
rect 185 505 200 575
rect 220 505 235 575
rect 185 490 235 505
rect -50 300 0 315
rect -50 230 -35 300
rect -15 230 0 300
rect -50 215 0 230
rect 15 300 65 315
rect 15 230 30 300
rect 50 230 65 300
rect 15 215 65 230
rect 80 300 130 315
rect 80 230 95 300
rect 115 230 130 300
rect 80 215 130 230
rect 145 215 170 315
rect 185 300 235 315
rect 185 230 200 300
rect 220 230 235 300
rect 185 215 235 230
<< ndiffc >>
rect -35 75 -15 145
rect 70 75 90 145
rect 135 75 155 145
rect 200 75 220 145
rect -35 -200 -15 -130
rect 70 -200 90 -130
rect 135 -200 155 -130
rect 200 -200 220 -130
<< pdiffc >>
rect -35 505 -15 575
rect 30 505 50 575
rect 95 505 115 575
rect 200 505 220 575
rect -35 230 -15 300
rect 30 230 50 300
rect 95 230 115 300
rect 200 230 220 300
<< psubdiff >>
rect -65 5 -15 20
rect -65 -65 -50 5
rect -30 -65 -15 5
rect -65 -80 -15 -65
<< nsubdiff >>
rect -60 440 -10 455
rect -60 370 -45 440
rect -25 370 -10 440
rect -60 355 -10 370
<< psubdiffcont >>
rect -50 -65 -30 5
<< nsubdiffcont >>
rect -45 370 -25 440
<< poly >>
rect 170 635 210 645
rect 170 615 180 635
rect 200 615 210 635
rect 170 605 210 615
rect 0 590 15 605
rect 65 590 80 605
rect 130 590 145 605
rect 170 590 185 605
rect 0 315 15 490
rect 65 475 80 490
rect 65 465 105 475
rect 65 445 75 465
rect 95 445 105 465
rect 65 435 105 445
rect 40 400 80 410
rect 40 380 50 400
rect 70 380 80 400
rect 40 370 80 380
rect 65 315 80 370
rect 130 315 145 490
rect 170 475 185 490
rect 190 420 230 430
rect 190 400 200 420
rect 220 400 230 420
rect 190 390 230 400
rect 190 340 210 390
rect 170 325 210 340
rect 170 315 185 325
rect 0 160 15 215
rect 65 200 80 215
rect 130 200 145 215
rect 40 185 80 200
rect 105 185 145 200
rect 40 160 55 185
rect 105 160 120 185
rect 170 160 185 215
rect 0 -115 15 60
rect 40 -10 55 60
rect 40 -20 80 -10
rect 40 -40 50 -20
rect 70 -40 80 -20
rect 40 -50 80 -40
rect 40 -115 55 -100
rect 105 -115 120 60
rect 170 5 185 60
rect 145 -5 185 5
rect 145 -25 155 -5
rect 175 -25 185 -5
rect 145 -35 185 -25
rect 170 -70 210 -60
rect 170 -90 180 -70
rect 200 -90 210 -70
rect 170 -100 210 -90
rect 170 -115 185 -100
rect 0 -270 15 -215
rect 40 -230 55 -215
rect 40 -240 80 -230
rect 40 -260 50 -240
rect 70 -260 80 -240
rect 40 -270 80 -260
rect 105 -270 120 -215
rect 170 -230 185 -215
rect -25 -280 15 -270
rect -25 -300 -15 -280
rect 5 -300 15 -280
rect -25 -310 15 -300
rect 105 -280 145 -270
rect 105 -300 115 -280
rect 135 -300 145 -280
rect 105 -310 145 -300
<< polycont >>
rect 180 615 200 635
rect 75 445 95 465
rect 50 380 70 400
rect 200 400 220 420
rect 50 -40 70 -20
rect 155 -25 175 -5
rect 180 -90 200 -70
rect 50 -260 70 -240
rect -15 -300 5 -280
rect 115 -300 135 -280
<< locali >>
rect 170 635 210 645
rect 170 625 180 635
rect 145 615 180 625
rect 200 615 210 635
rect 145 605 210 615
rect -45 575 -5 585
rect -45 515 -35 575
rect -85 505 -35 515
rect -15 505 -5 575
rect -85 495 -5 505
rect 20 575 60 585
rect 20 505 30 575
rect 50 505 60 575
rect 20 495 60 505
rect 85 575 125 585
rect 85 505 95 575
rect 115 505 125 575
rect 85 495 125 505
rect -55 440 -15 450
rect -55 370 -45 440
rect -25 370 -15 440
rect 20 410 40 495
rect 65 465 105 475
rect 65 445 75 465
rect 95 455 105 465
rect 95 445 120 455
rect 65 435 120 445
rect 20 400 80 410
rect 20 390 50 400
rect 40 380 50 390
rect 70 380 80 400
rect 40 370 80 380
rect -55 360 -15 370
rect 100 350 120 435
rect 40 330 120 350
rect 40 310 60 330
rect 145 310 165 605
rect 190 575 230 585
rect 190 505 200 575
rect 220 515 230 575
rect 220 505 255 515
rect 190 495 255 505
rect 210 430 230 495
rect 190 420 230 430
rect 190 400 200 420
rect 220 400 230 420
rect 190 390 230 400
rect -85 300 -5 310
rect -85 290 -35 300
rect -45 230 -35 290
rect -15 230 -5 300
rect -45 220 -5 230
rect 20 300 60 310
rect 20 230 30 300
rect 50 230 60 300
rect 20 220 60 230
rect 85 300 125 310
rect 85 230 95 300
rect 115 230 125 300
rect 145 300 255 310
rect 145 290 200 300
rect 85 220 125 230
rect 190 230 200 290
rect 220 290 255 300
rect 220 230 230 290
rect 190 220 230 230
rect 40 195 60 220
rect 190 195 210 220
rect 40 175 80 195
rect 60 155 80 175
rect 145 175 210 195
rect 145 155 165 175
rect -45 145 -5 155
rect -45 75 -35 145
rect -15 75 -5 145
rect 60 145 100 155
rect 60 85 70 145
rect -45 65 -5 75
rect 15 75 70 85
rect 90 75 100 145
rect 15 65 100 75
rect 125 145 165 155
rect 125 75 135 145
rect 155 75 165 145
rect 125 65 165 75
rect 190 145 230 155
rect 190 75 200 145
rect 220 75 230 145
rect 190 65 230 75
rect 15 45 35 65
rect 0 25 35 45
rect 145 45 165 65
rect 145 25 225 45
rect -60 5 -20 15
rect -60 -65 -50 5
rect -30 -65 -20 5
rect -60 -75 -20 -65
rect 0 -80 20 25
rect 145 -5 185 5
rect 40 -20 80 -10
rect 145 -15 155 -5
rect 40 -40 50 -20
rect 70 -40 80 -20
rect 40 -50 80 -40
rect 0 -100 35 -80
rect -45 -130 -5 -120
rect -45 -200 -35 -130
rect -15 -200 -5 -130
rect -45 -210 -5 -200
rect 15 -230 35 -100
rect 60 -120 80 -50
rect 125 -25 155 -15
rect 175 -25 185 -5
rect 125 -35 185 -25
rect 125 -120 145 -35
rect 205 -60 225 25
rect 170 -70 225 -60
rect 170 -90 180 -70
rect 200 -80 225 -70
rect 200 -90 210 -80
rect 170 -100 210 -90
rect 60 -130 100 -120
rect 60 -200 70 -130
rect 90 -200 100 -130
rect 60 -210 100 -200
rect 125 -130 165 -120
rect 125 -200 135 -130
rect 155 -200 165 -130
rect 125 -210 165 -200
rect 190 -130 230 -120
rect 190 -200 200 -130
rect 220 -200 230 -130
rect 190 -210 230 -200
rect 15 -240 80 -230
rect 15 -250 50 -240
rect 40 -260 50 -250
rect 70 -260 80 -240
rect 40 -270 80 -260
rect -25 -280 15 -270
rect -25 -300 -15 -280
rect 5 -300 15 -280
rect -25 -310 15 -300
rect 105 -280 145 -270
rect 105 -300 115 -280
rect 135 -300 145 -280
rect 105 -310 145 -300
<< viali >>
rect 95 505 115 575
rect -45 370 -25 440
rect 95 230 115 300
rect -35 75 -15 145
rect 200 75 220 145
rect -50 -65 -30 5
rect -35 -200 -15 -130
rect 200 -200 220 -130
rect -15 -300 5 -280
rect 115 -300 135 -280
<< metal1 >>
rect -85 575 255 590
rect -85 505 95 575
rect 115 505 255 575
rect -85 440 255 505
rect -85 370 -45 440
rect -25 370 255 440
rect -85 300 255 370
rect -85 230 95 300
rect 115 230 255 300
rect -85 215 255 230
rect -85 145 255 160
rect -85 75 -35 145
rect -15 75 200 145
rect 220 75 255 145
rect -85 5 255 75
rect -85 -65 -50 5
rect -30 -65 255 5
rect -85 -130 255 -65
rect -85 -200 -35 -130
rect -15 -200 200 -130
rect 220 -200 255 -130
rect -85 -215 255 -200
rect -85 -280 255 -270
rect -85 -300 -15 -280
rect 5 -300 115 -280
rect 135 -300 255 -280
rect -85 -310 255 -300
<< labels >>
rlabel metal1 -85 -40 -85 -40 7 VN
rlabel metal1 -85 400 -85 400 7 VP
rlabel locali -85 300 -85 300 7 D
rlabel locali -85 505 -85 505 7 nD
rlabel locali 255 300 255 300 3 Q
rlabel locali 255 505 255 505 3 nQ
rlabel metal1 -85 -290 -85 -290 7 CLK
<< end >>
