magic
tech sky130A
timestamp 1615439024
<< nwell >>
rect -520 1225 670 4085
<< nmos >>
rect -400 440 -350 1040
rect -300 440 -250 1040
rect -200 440 -150 1040
rect -100 440 -50 1040
rect 0 440 50 1040
rect 100 440 150 1040
rect 200 440 250 1040
rect 300 440 350 1040
rect 400 440 450 1040
rect 500 440 550 1040
<< pmos >>
rect -400 3465 -350 4065
rect -300 3465 -250 4065
rect -200 3465 -150 4065
rect -100 3465 -50 4065
rect 0 3465 50 4065
rect 100 3465 150 4065
rect 200 3465 250 4065
rect 300 3465 350 4065
rect 400 3465 450 4065
rect 500 3465 550 4065
rect -400 2090 -350 3290
rect -300 2090 -250 3290
rect -200 2090 -150 3290
rect -100 2090 -50 3290
rect 0 2090 50 3290
rect 100 2090 150 3290
rect 200 2090 250 3290
rect 300 2090 350 3290
rect 400 2090 450 3290
rect 500 2090 550 3290
rect -400 1245 -350 1845
rect -300 1245 -250 1845
rect -200 1245 -150 1845
rect -100 1245 -50 1845
rect 0 1245 50 1845
rect 100 1245 150 1845
rect 200 1245 250 1845
rect 300 1245 350 1845
rect 400 1245 450 1845
rect 500 1245 550 1845
<< ndiff >>
rect -450 1025 -400 1040
rect -450 455 -435 1025
rect -415 455 -400 1025
rect -450 440 -400 455
rect -350 1025 -300 1040
rect -350 455 -335 1025
rect -315 455 -300 1025
rect -350 440 -300 455
rect -250 1025 -200 1040
rect -250 455 -235 1025
rect -215 455 -200 1025
rect -250 440 -200 455
rect -150 1025 -100 1040
rect -150 455 -135 1025
rect -115 455 -100 1025
rect -150 440 -100 455
rect -50 1025 0 1040
rect -50 455 -35 1025
rect -15 455 0 1025
rect -50 440 0 455
rect 50 1025 100 1040
rect 50 455 65 1025
rect 85 455 100 1025
rect 50 440 100 455
rect 150 1025 200 1040
rect 150 455 165 1025
rect 185 455 200 1025
rect 150 440 200 455
rect 250 1025 300 1040
rect 250 455 265 1025
rect 285 455 300 1025
rect 250 440 300 455
rect 350 1025 400 1040
rect 350 455 365 1025
rect 385 455 400 1025
rect 350 440 400 455
rect 450 1025 500 1040
rect 450 455 465 1025
rect 485 455 500 1025
rect 450 440 500 455
rect 550 1025 600 1040
rect 550 455 565 1025
rect 585 455 600 1025
rect 550 440 600 455
<< pdiff >>
rect -450 4050 -400 4065
rect -450 3480 -435 4050
rect -415 3480 -400 4050
rect -450 3465 -400 3480
rect -350 4050 -300 4065
rect -350 3480 -335 4050
rect -315 3480 -300 4050
rect -350 3465 -300 3480
rect -250 4050 -200 4065
rect -250 3480 -235 4050
rect -215 3480 -200 4050
rect -250 3465 -200 3480
rect -150 4050 -100 4065
rect -150 3480 -135 4050
rect -115 3480 -100 4050
rect -150 3465 -100 3480
rect -50 4050 0 4065
rect -50 3480 -35 4050
rect -15 3480 0 4050
rect -50 3465 0 3480
rect 50 4050 100 4065
rect 50 3480 65 4050
rect 85 3480 100 4050
rect 50 3465 100 3480
rect 150 4050 200 4065
rect 150 3480 165 4050
rect 185 3480 200 4050
rect 150 3465 200 3480
rect 250 4050 300 4065
rect 250 3480 265 4050
rect 285 3480 300 4050
rect 250 3465 300 3480
rect 350 4050 400 4065
rect 350 3480 365 4050
rect 385 3480 400 4050
rect 350 3465 400 3480
rect 450 4050 500 4065
rect 450 3480 465 4050
rect 485 3480 500 4050
rect 450 3465 500 3480
rect 550 4050 600 4065
rect 550 3480 565 4050
rect 585 3480 600 4050
rect 550 3465 600 3480
rect -450 3275 -400 3290
rect -450 2105 -435 3275
rect -415 2105 -400 3275
rect -450 2090 -400 2105
rect -350 3275 -300 3290
rect -350 2105 -335 3275
rect -315 2105 -300 3275
rect -350 2090 -300 2105
rect -250 3275 -200 3290
rect -250 2105 -235 3275
rect -215 2105 -200 3275
rect -250 2090 -200 2105
rect -150 3275 -100 3290
rect -150 2105 -135 3275
rect -115 2105 -100 3275
rect -150 2090 -100 2105
rect -50 3275 0 3290
rect -50 2105 -35 3275
rect -15 2105 0 3275
rect -50 2090 0 2105
rect 50 3275 100 3290
rect 50 2105 65 3275
rect 85 2105 100 3275
rect 50 2090 100 2105
rect 150 3275 200 3290
rect 150 2105 165 3275
rect 185 2105 200 3275
rect 150 2090 200 2105
rect 250 3275 300 3290
rect 250 2105 265 3275
rect 285 2105 300 3275
rect 250 2090 300 2105
rect 350 3275 400 3290
rect 350 2105 365 3275
rect 385 2105 400 3275
rect 350 2090 400 2105
rect 450 3275 500 3290
rect 450 2105 465 3275
rect 485 2105 500 3275
rect 450 2090 500 2105
rect 550 3275 600 3290
rect 550 2105 565 3275
rect 585 2105 600 3275
rect 550 2090 600 2105
rect -450 1830 -400 1845
rect -450 1260 -435 1830
rect -415 1260 -400 1830
rect -450 1245 -400 1260
rect -350 1830 -300 1845
rect -350 1260 -335 1830
rect -315 1260 -300 1830
rect -350 1245 -300 1260
rect -250 1830 -200 1845
rect -250 1260 -235 1830
rect -215 1260 -200 1830
rect -250 1245 -200 1260
rect -150 1830 -100 1845
rect -150 1260 -135 1830
rect -115 1260 -100 1830
rect -150 1245 -100 1260
rect -50 1830 0 1845
rect -50 1260 -35 1830
rect -15 1260 0 1830
rect -50 1245 0 1260
rect 50 1830 100 1845
rect 50 1260 65 1830
rect 85 1260 100 1830
rect 50 1245 100 1260
rect 150 1830 200 1845
rect 150 1260 165 1830
rect 185 1260 200 1830
rect 150 1245 200 1260
rect 250 1830 300 1845
rect 250 1260 265 1830
rect 285 1260 300 1830
rect 250 1245 300 1260
rect 350 1830 400 1845
rect 350 1260 365 1830
rect 385 1260 400 1830
rect 350 1245 400 1260
rect 450 1830 500 1845
rect 450 1260 465 1830
rect 485 1260 500 1830
rect 450 1245 500 1260
rect 550 1830 600 1845
rect 550 1260 565 1830
rect 585 1260 600 1830
rect 550 1245 600 1260
<< ndiffc >>
rect -435 455 -415 1025
rect -335 455 -315 1025
rect -235 455 -215 1025
rect -135 455 -115 1025
rect -35 455 -15 1025
rect 65 455 85 1025
rect 165 455 185 1025
rect 265 455 285 1025
rect 365 455 385 1025
rect 465 455 485 1025
rect 565 455 585 1025
<< pdiffc >>
rect -435 3480 -415 4050
rect -335 3480 -315 4050
rect -235 3480 -215 4050
rect -135 3480 -115 4050
rect -35 3480 -15 4050
rect 65 3480 85 4050
rect 165 3480 185 4050
rect 265 3480 285 4050
rect 365 3480 385 4050
rect 465 3480 485 4050
rect 565 3480 585 4050
rect -435 2105 -415 3275
rect -335 2105 -315 3275
rect -235 2105 -215 3275
rect -135 2105 -115 3275
rect -35 2105 -15 3275
rect 65 2105 85 3275
rect 165 2105 185 3275
rect 265 2105 285 3275
rect 365 2105 385 3275
rect 465 2105 485 3275
rect 565 2105 585 3275
rect -435 1260 -415 1830
rect -335 1260 -315 1830
rect -235 1260 -215 1830
rect -135 1260 -115 1830
rect -35 1260 -15 1830
rect 65 1260 85 1830
rect 165 1260 185 1830
rect 265 1260 285 1830
rect 365 1260 385 1830
rect 465 1260 485 1830
rect 565 1260 585 1830
<< psubdiff >>
rect -500 1025 -450 1040
rect -500 455 -485 1025
rect -465 455 -450 1025
rect -500 440 -450 455
rect 600 1025 650 1040
rect 600 455 615 1025
rect 635 455 650 1025
rect 600 440 650 455
<< nsubdiff >>
rect -500 4050 -450 4065
rect -500 3480 -485 4050
rect -465 3480 -450 4050
rect -500 3465 -450 3480
rect 600 4050 650 4065
rect 600 3480 615 4050
rect 635 3480 650 4050
rect 600 3465 650 3480
rect -500 3275 -450 3290
rect -500 2105 -485 3275
rect -465 2105 -450 3275
rect -500 2090 -450 2105
rect 600 3275 650 3290
rect 600 2105 615 3275
rect 635 2105 650 3275
rect 600 2090 650 2105
rect -500 1830 -450 1845
rect -500 1260 -485 1830
rect -465 1260 -450 1830
rect -500 1245 -450 1260
rect 600 1830 650 1845
rect 600 1260 615 1830
rect 635 1260 650 1830
rect 600 1245 650 1260
<< psubdiffcont >>
rect -485 455 -465 1025
rect 615 455 635 1025
<< nsubdiffcont >>
rect -485 3480 -465 4050
rect 615 3480 635 4050
rect -485 2105 -465 3275
rect 615 2105 635 3275
rect -485 1260 -465 1830
rect 615 1260 635 1830
<< poly >>
rect -500 4150 450 4200
rect -450 4110 -350 4125
rect -450 4090 -435 4110
rect -415 4090 -350 4110
rect -450 4075 -350 4090
rect -400 4065 -350 4075
rect -300 4065 -250 4150
rect -200 4065 -150 4150
rect -100 4065 -50 4150
rect 0 4065 50 4150
rect 100 4065 150 4150
rect 200 4065 250 4150
rect 300 4065 350 4150
rect 400 4065 450 4150
rect 500 4110 600 4125
rect 500 4090 565 4110
rect 585 4090 600 4110
rect 500 4075 600 4090
rect 500 4065 550 4075
rect -400 3450 -350 3465
rect -300 3450 -250 3465
rect -200 3450 -150 3465
rect -100 3450 -50 3465
rect 0 3450 50 3465
rect 100 3450 150 3465
rect 200 3450 250 3465
rect 300 3450 350 3465
rect 400 3450 450 3465
rect 500 3450 550 3465
rect -500 3375 450 3425
rect -450 3335 -350 3350
rect -450 3315 -435 3335
rect -415 3315 -350 3335
rect -450 3300 -350 3315
rect -400 3290 -350 3300
rect -300 3290 -250 3375
rect -200 3290 -150 3375
rect -100 3290 -50 3305
rect 0 3290 50 3305
rect 100 3290 150 3305
rect 200 3290 250 3305
rect 300 3290 350 3375
rect 400 3290 450 3375
rect 500 3335 600 3350
rect 500 3315 565 3335
rect 585 3315 600 3335
rect 500 3300 600 3315
rect 500 3290 550 3300
rect -400 2075 -350 2090
rect -300 2075 -250 2090
rect -200 2075 -150 2090
rect -100 2050 -50 2090
rect 0 2050 50 2090
rect 100 2050 150 2090
rect 200 2050 250 2090
rect 300 2075 350 2090
rect 400 2075 450 2090
rect 500 2075 550 2090
rect -500 2005 250 2050
rect -500 1930 450 1980
rect -450 1890 -350 1905
rect -450 1870 -435 1890
rect -415 1870 -350 1890
rect -450 1855 -350 1870
rect -400 1845 -350 1855
rect -300 1845 -250 1930
rect -200 1845 -150 1860
rect -100 1845 -50 1860
rect 0 1845 50 1930
rect 100 1845 150 1930
rect 200 1845 250 1860
rect 300 1845 350 1860
rect 400 1845 450 1930
rect 500 1890 600 1905
rect 500 1870 565 1890
rect 585 1870 600 1890
rect 500 1855 600 1870
rect 500 1845 550 1855
rect -400 1230 -350 1245
rect -300 1230 -250 1245
rect -200 1205 -150 1245
rect -100 1205 -50 1245
rect 0 1230 50 1245
rect 100 1230 150 1245
rect 200 1205 250 1245
rect 300 1205 350 1245
rect 400 1230 450 1245
rect 500 1230 550 1245
rect -200 1190 350 1205
rect -200 1170 65 1190
rect 85 1170 350 1190
rect -200 1155 350 1170
rect -500 1080 350 1130
rect -400 1040 -350 1055
rect -300 1040 -250 1055
rect -200 1040 -150 1080
rect -100 1040 -50 1080
rect 0 1040 50 1055
rect 100 1040 150 1055
rect 200 1040 250 1080
rect 300 1040 350 1080
rect 400 1040 450 1055
rect 500 1040 550 1055
rect -400 430 -350 440
rect -450 415 -350 430
rect -450 395 -435 415
rect -415 395 -350 415
rect -450 380 -350 395
rect -300 355 -250 440
rect -200 425 -150 440
rect -100 425 -50 440
rect 0 355 50 440
rect 100 355 150 440
rect 200 425 250 440
rect 300 425 350 440
rect 400 355 450 440
rect 500 430 550 440
rect 500 415 600 430
rect 500 395 565 415
rect 585 395 600 415
rect 500 380 600 395
rect -500 305 450 355
<< polycont >>
rect -435 4090 -415 4110
rect 565 4090 585 4110
rect -435 3315 -415 3335
rect 565 3315 585 3335
rect -435 1870 -415 1890
rect 565 1870 585 1890
rect 65 1170 85 1190
rect -435 395 -415 415
rect 565 395 585 415
<< locali >>
rect -445 4110 -405 4120
rect -445 4090 -435 4110
rect -415 4090 -405 4110
rect -445 4060 -405 4090
rect 555 4110 595 4120
rect 555 4090 565 4110
rect 585 4090 595 4110
rect 555 4060 595 4090
rect -495 4050 -405 4060
rect -495 3480 -485 4050
rect -465 3480 -435 4050
rect -415 3480 -405 4050
rect -495 3470 -405 3480
rect -345 4050 -305 4060
rect -345 3480 -335 4050
rect -315 3480 -305 4050
rect -345 3470 -305 3480
rect -245 4050 -205 4060
rect -245 3480 -235 4050
rect -215 3480 -205 4050
rect -245 3470 -205 3480
rect -145 4050 -105 4060
rect -145 3480 -135 4050
rect -115 3480 -105 4050
rect -145 3445 -105 3480
rect -45 4050 -5 4060
rect -45 3480 -35 4050
rect -15 3480 -5 4050
rect -45 3470 -5 3480
rect 55 4050 95 4060
rect 55 3480 65 4050
rect 85 3480 95 4050
rect 55 3470 95 3480
rect 155 4050 195 4060
rect 155 3480 165 4050
rect 185 3480 195 4050
rect 155 3470 195 3480
rect 255 4050 295 4060
rect 255 3480 265 4050
rect 285 3480 295 4050
rect 255 3445 295 3480
rect 355 4050 395 4060
rect 355 3480 365 4050
rect 385 3480 395 4050
rect 355 3470 395 3480
rect 455 4050 495 4060
rect 455 3480 465 4050
rect 485 3480 495 4050
rect 455 3470 495 3480
rect 555 4050 645 4060
rect 555 3480 565 4050
rect 585 3480 615 4050
rect 635 3480 645 4050
rect 555 3470 645 3480
rect -145 3405 295 3445
rect -445 3335 -405 3345
rect -445 3315 -435 3335
rect -415 3315 -405 3335
rect -445 3285 -405 3315
rect -495 3275 -405 3285
rect -495 2105 -485 3275
rect -465 2105 -435 3275
rect -415 2105 -405 3275
rect -495 2095 -405 2105
rect -345 3275 -305 3285
rect -345 2105 -335 3275
rect -315 2105 -305 3275
rect -345 2095 -305 2105
rect -245 3275 -205 3285
rect -245 2105 -235 3275
rect -215 2105 -205 3275
rect -245 2095 -205 2105
rect -145 3275 -105 3405
rect -145 2105 -135 3275
rect -115 2105 -105 3275
rect -145 2095 -105 2105
rect -45 3275 -5 3285
rect -45 2105 -35 3275
rect -15 2105 -5 3275
rect -45 2095 -5 2105
rect 55 3275 95 3285
rect 55 2105 65 3275
rect 85 2105 95 3275
rect 55 2095 95 2105
rect 155 3275 195 3285
rect 155 2105 165 3275
rect 185 2105 195 3275
rect 155 2095 195 2105
rect 255 3275 295 3405
rect 555 3335 595 3345
rect 555 3315 565 3335
rect 585 3315 595 3335
rect 555 3285 595 3315
rect 255 2105 265 3275
rect 285 2105 295 3275
rect 255 2095 295 2105
rect 355 3275 395 3285
rect 355 2105 365 3275
rect 385 2105 395 3275
rect 355 2095 395 2105
rect 455 3275 495 3285
rect 455 2105 465 3275
rect 485 2105 495 3275
rect 455 2095 495 2105
rect 555 3275 645 3285
rect 555 2105 565 3275
rect 585 2105 615 3275
rect 635 2105 645 3275
rect 555 2095 645 2105
rect -445 1890 -405 1900
rect -445 1870 -435 1890
rect -415 1870 -405 1890
rect -445 1840 -405 1870
rect -495 1830 -405 1840
rect -495 1260 -485 1830
rect -465 1260 -435 1830
rect -415 1260 -405 1830
rect -495 1250 -405 1260
rect -345 1860 495 1900
rect -345 1830 -305 1860
rect -345 1260 -335 1830
rect -315 1260 -305 1830
rect -495 1025 -405 1035
rect -495 455 -485 1025
rect -465 455 -435 1025
rect -415 455 -405 1025
rect -495 445 -405 455
rect -445 415 -405 445
rect -445 395 -435 415
rect -415 395 -405 415
rect -445 385 -405 395
rect -345 1025 -305 1260
rect -245 1830 -205 1840
rect -245 1260 -235 1830
rect -215 1260 -205 1830
rect -245 1250 -205 1260
rect -145 1830 -105 1840
rect -145 1260 -135 1830
rect -115 1260 -105 1830
rect -145 1250 -105 1260
rect -45 1830 -5 1840
rect -45 1260 -35 1830
rect -15 1260 -5 1830
rect -45 1250 -5 1260
rect 55 1830 95 1840
rect 55 1260 65 1830
rect 85 1260 95 1830
rect 55 1190 95 1260
rect 155 1830 195 1840
rect 155 1260 165 1830
rect 185 1260 195 1830
rect 155 1250 195 1260
rect 255 1830 295 1840
rect 255 1260 265 1830
rect 285 1260 295 1830
rect 255 1250 295 1260
rect 355 1830 395 1840
rect 355 1260 365 1830
rect 385 1260 395 1830
rect 355 1250 395 1260
rect 455 1830 495 1860
rect 455 1260 465 1830
rect 485 1260 495 1830
rect 55 1170 65 1190
rect 85 1170 95 1190
rect -345 455 -335 1025
rect -315 455 -305 1025
rect -345 365 -305 455
rect -245 1025 -205 1035
rect -245 455 -235 1025
rect -215 455 -205 1025
rect -245 425 -205 455
rect -145 1025 -105 1035
rect -145 455 -135 1025
rect -115 455 -105 1025
rect -145 445 -105 455
rect -45 1025 -5 1035
rect -45 455 -35 1025
rect -15 455 -5 1025
rect -45 445 -5 455
rect 55 1025 95 1170
rect 455 1165 495 1260
rect 555 1890 595 1900
rect 555 1870 565 1890
rect 585 1870 595 1890
rect 555 1840 595 1870
rect 555 1830 645 1840
rect 555 1260 565 1830
rect 585 1260 615 1830
rect 635 1260 645 1830
rect 555 1250 645 1260
rect 455 1125 650 1165
rect 55 455 65 1025
rect 85 455 95 1025
rect 55 445 95 455
rect 155 1025 195 1035
rect 155 455 165 1025
rect 185 455 195 1025
rect 155 445 195 455
rect 255 1025 295 1035
rect 255 455 265 1025
rect 285 455 295 1025
rect 255 445 295 455
rect 355 1025 395 1035
rect 355 455 365 1025
rect 385 455 395 1025
rect 355 425 395 455
rect -245 385 395 425
rect 455 1025 495 1125
rect 455 455 465 1025
rect 485 455 495 1025
rect 455 365 495 455
rect 555 1025 645 1035
rect 555 455 565 1025
rect 585 455 615 1025
rect 635 455 645 1025
rect 555 445 645 455
rect 555 415 595 445
rect 555 395 565 415
rect 585 395 595 415
rect 555 385 595 395
rect -345 325 495 365
<< viali >>
rect -485 3480 -465 4050
rect -435 3480 -415 4050
rect -335 3480 -315 4050
rect 65 3480 85 4050
rect 465 3480 485 4050
rect 565 3480 585 4050
rect 615 3480 635 4050
rect -485 2105 -465 3275
rect -435 2105 -415 3275
rect -335 2105 -315 3275
rect 65 2105 85 3275
rect 465 2105 485 3275
rect 565 2105 585 3275
rect 615 2105 635 3275
rect -485 1260 -465 1830
rect -435 1260 -415 1830
rect -485 455 -465 1025
rect -435 455 -415 1025
rect -135 1260 -115 1830
rect 265 1260 285 1830
rect -235 455 -215 1025
rect -135 455 -115 1025
rect -35 455 -15 1025
rect 565 1260 585 1830
rect 615 1260 635 1830
rect 165 455 185 1025
rect 265 455 285 1025
rect 365 455 385 1025
rect 565 455 585 1025
rect 615 455 635 1025
<< metal1 >>
rect -500 4100 650 4250
rect -495 4050 -405 4100
rect -495 3480 -485 4050
rect -465 3480 -435 4050
rect -415 3480 -405 4050
rect -495 3275 -405 3480
rect -345 4050 -305 4100
rect -345 3480 -335 4050
rect -315 3480 -305 4050
rect -345 3470 -305 3480
rect -495 2105 -485 3275
rect -465 2105 -435 3275
rect -415 2105 -405 3275
rect -495 1830 -405 2105
rect -495 1260 -485 1830
rect -465 1260 -435 1830
rect -415 1260 -405 1830
rect -495 1250 -405 1260
rect -345 3275 -305 3285
rect -345 2105 -335 3275
rect -315 2105 -305 3275
rect -345 1165 -305 2105
rect -145 1830 -105 4100
rect 55 4050 95 4100
rect 55 3480 65 4050
rect 85 3480 95 4050
rect 55 3470 95 3480
rect 55 3275 95 3285
rect 55 2105 65 3275
rect 85 2105 95 3275
rect 55 2020 95 2105
rect -145 1260 -135 1830
rect -115 1260 -105 1830
rect -145 1250 -105 1260
rect -45 1980 195 2020
rect -345 1125 -205 1165
rect -495 1025 -405 1035
rect -495 455 -485 1025
rect -465 455 -435 1025
rect -415 455 -405 1025
rect -495 405 -405 455
rect -245 1025 -205 1125
rect -245 455 -235 1025
rect -215 455 -205 1025
rect -245 445 -205 455
rect -145 1025 -105 1035
rect -145 455 -135 1025
rect -115 455 -105 1025
rect -145 405 -105 455
rect -45 1025 -5 1980
rect -45 455 -35 1025
rect -15 455 -5 1025
rect -45 445 -5 455
rect 155 1025 195 1980
rect 255 1830 295 4100
rect 455 4050 495 4100
rect 455 3480 465 4050
rect 485 3480 495 4050
rect 455 3470 495 3480
rect 555 4050 645 4100
rect 555 3480 565 4050
rect 585 3480 615 4050
rect 635 3480 645 4050
rect 255 1260 265 1830
rect 285 1260 295 1830
rect 255 1250 295 1260
rect 455 3275 495 3285
rect 455 2105 465 3275
rect 485 2105 495 3275
rect 455 1165 495 2105
rect 555 3275 645 3480
rect 555 2105 565 3275
rect 585 2105 615 3275
rect 635 2105 645 3275
rect 555 1830 645 2105
rect 555 1260 565 1830
rect 585 1260 615 1830
rect 635 1260 645 1830
rect 555 1250 645 1260
rect 355 1125 495 1165
rect 155 455 165 1025
rect 185 455 195 1025
rect 155 445 195 455
rect 255 1025 295 1035
rect 255 455 265 1025
rect 285 455 295 1025
rect 255 405 295 455
rect 355 1025 395 1125
rect 355 455 365 1025
rect 385 455 395 1025
rect 355 445 395 455
rect 555 1025 645 1035
rect 555 455 565 1025
rect 585 455 615 1025
rect 635 455 645 1025
rect 555 405 645 455
rect -500 255 650 405
<< labels >>
rlabel metal1 -500 4170 -500 4170 3 VDD
rlabel poly -500 4175 -500 4175 7 Vbp
rlabel poly -500 3400 -500 3400 7 V2
rlabel pdiff -225 3465 -225 3465 5 net7
rlabel locali -125 4060 -125 4060 1 net8
rlabel poly -500 1955 -500 1955 7 Vcp
rlabel poly -500 330 -500 330 7 Vcn
rlabel metal1 -500 290 -500 290 3 GND
rlabel poly -500 2025 -500 2025 7 V1
rlabel poly -500 1100 -500 1100 7 Vbn
rlabel locali 375 3470 375 3470 5 net11
rlabel pdiff 175 2090 175 2090 5 net14
rlabel pdiff -25 2090 -25 2090 5 net13
rlabel pdiff -225 2090 -225 2090 5 net15
rlabel pdiff 375 2090 375 2090 5 net16
rlabel pdiff 375 1245 375 1245 5 net6
<< end >>
