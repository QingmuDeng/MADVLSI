magic
tech sky130A
timestamp 1612841356
<< nwell >>
rect -145 140 125 280
<< nmos >>
rect 0 0 15 100
rect 40 0 55 100
<< pmos >>
rect -25 160 -10 260
rect 40 160 55 260
<< ndiff >>
rect -50 85 0 100
rect -50 15 -35 85
rect -15 15 0 85
rect -50 0 0 15
rect 15 0 40 100
rect 55 85 105 100
rect 55 15 70 85
rect 90 15 105 85
rect 55 0 105 15
<< pdiff >>
rect -75 245 -25 260
rect -75 175 -60 245
rect -40 175 -25 245
rect -75 160 -25 175
rect -10 245 40 260
rect -10 175 5 245
rect 25 175 40 245
rect -10 160 40 175
rect 55 245 105 260
rect 55 175 70 245
rect 90 175 105 245
rect 55 160 105 175
<< ndiffc >>
rect -35 15 -15 85
rect 70 15 90 85
<< pdiffc >>
rect -60 175 -40 245
rect 5 175 25 245
rect 70 175 90 245
<< psubdiff >>
rect -130 85 -80 100
rect -130 15 -115 85
rect -95 15 -80 85
rect -130 0 -80 15
<< nsubdiff >>
rect -125 245 -75 260
rect -125 175 -110 245
rect -90 175 -75 245
rect -125 160 -75 175
<< psubdiffcont >>
rect -115 15 -95 85
<< nsubdiffcont >>
rect -110 175 -90 245
<< poly >>
rect 15 305 55 315
rect 15 285 25 305
rect 45 285 55 305
rect 15 275 55 285
rect -25 260 -10 275
rect 40 260 55 275
rect -25 135 -10 160
rect -25 120 15 135
rect 0 100 15 120
rect 40 100 55 160
rect 0 -15 15 0
rect 40 -15 55 0
rect -25 -25 15 -15
rect -25 -45 -15 -25
rect 5 -45 15 -25
rect -25 -55 15 -45
<< polycont >>
rect 25 285 45 305
rect -15 -45 5 -25
<< locali >>
rect 15 305 55 315
rect 15 295 25 305
rect -145 285 25 295
rect 45 285 55 305
rect -145 275 55 285
rect -120 245 -30 255
rect -120 175 -110 245
rect -90 175 -60 245
rect -40 175 -30 245
rect -120 165 -30 175
rect -5 245 35 255
rect -5 175 5 245
rect 25 175 35 245
rect -5 165 35 175
rect 60 245 100 255
rect 60 175 70 245
rect 90 175 100 245
rect 60 165 100 175
rect 15 140 35 165
rect 15 120 100 140
rect 80 95 100 120
rect -125 85 -85 95
rect -125 15 -115 85
rect -95 15 -85 85
rect -125 5 -85 15
rect -45 85 -5 95
rect -45 15 -35 85
rect -15 15 -5 85
rect -45 5 -5 15
rect 60 85 100 95
rect 60 15 70 85
rect 90 15 100 85
rect 60 5 100 15
rect 80 -15 100 5
rect -145 -25 15 -15
rect -145 -35 -15 -25
rect -25 -45 -15 -35
rect 5 -45 15 -25
rect 80 -35 125 -15
rect -25 -55 15 -45
<< end >>
