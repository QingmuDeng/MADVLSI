magic
tech sky130A
timestamp 1615756184
<< nwell >>
rect -520 1220 670 4085
<< nmos >>
rect -400 435 -350 1035
rect -300 435 -250 1035
rect -200 435 -150 1035
rect -100 435 -50 1035
rect 0 435 50 1035
rect 100 435 150 1035
rect 200 435 250 1035
rect 300 435 350 1035
rect 400 435 450 1035
rect 500 435 550 1035
<< pmos >>
rect -400 3465 -350 4065
rect -300 3465 -250 4065
rect -200 3465 -150 4065
rect -100 3465 -50 4065
rect 0 3465 50 4065
rect 100 3465 150 4065
rect 200 3465 250 4065
rect 300 3465 350 4065
rect 400 3465 450 4065
rect 500 3465 550 4065
rect -400 2090 -350 3290
rect -300 2090 -250 3290
rect -200 2090 -150 3290
rect -100 2090 -50 3290
rect 0 2090 50 3290
rect 100 2090 150 3290
rect 200 2090 250 3290
rect 300 2090 350 3290
rect 400 2090 450 3290
rect 500 2090 550 3290
rect -400 1240 -350 1840
rect -300 1240 -250 1840
rect -200 1240 -150 1840
rect -100 1240 -50 1840
rect 0 1240 50 1840
rect 100 1240 150 1840
rect 200 1240 250 1840
rect 300 1240 350 1840
rect 400 1240 450 1840
rect 500 1240 550 1840
<< ndiff >>
rect -450 1020 -400 1035
rect -450 450 -435 1020
rect -415 450 -400 1020
rect -450 435 -400 450
rect -350 1020 -300 1035
rect -350 450 -335 1020
rect -315 450 -300 1020
rect -350 435 -300 450
rect -250 1020 -200 1035
rect -250 450 -235 1020
rect -215 450 -200 1020
rect -250 435 -200 450
rect -150 1020 -100 1035
rect -150 450 -135 1020
rect -115 450 -100 1020
rect -150 435 -100 450
rect -50 1020 0 1035
rect -50 450 -35 1020
rect -15 450 0 1020
rect -50 435 0 450
rect 50 1020 100 1035
rect 50 450 65 1020
rect 85 450 100 1020
rect 50 435 100 450
rect 150 1020 200 1035
rect 150 450 165 1020
rect 185 450 200 1020
rect 150 435 200 450
rect 250 1020 300 1035
rect 250 450 265 1020
rect 285 450 300 1020
rect 250 435 300 450
rect 350 1020 400 1035
rect 350 450 365 1020
rect 385 450 400 1020
rect 350 435 400 450
rect 450 1020 500 1035
rect 450 450 465 1020
rect 485 450 500 1020
rect 450 435 500 450
rect 550 1020 600 1035
rect 550 450 565 1020
rect 585 450 600 1020
rect 550 435 600 450
<< pdiff >>
rect -450 4050 -400 4065
rect -450 3480 -435 4050
rect -415 3480 -400 4050
rect -450 3465 -400 3480
rect -350 4050 -300 4065
rect -350 3480 -335 4050
rect -315 3480 -300 4050
rect -350 3465 -300 3480
rect -250 4050 -200 4065
rect -250 3480 -235 4050
rect -215 3480 -200 4050
rect -250 3465 -200 3480
rect -150 4050 -100 4065
rect -150 3480 -135 4050
rect -115 3480 -100 4050
rect -150 3465 -100 3480
rect -50 4050 0 4065
rect -50 3480 -35 4050
rect -15 3480 0 4050
rect -50 3465 0 3480
rect 50 4050 100 4065
rect 50 3480 65 4050
rect 85 3480 100 4050
rect 50 3465 100 3480
rect 150 4050 200 4065
rect 150 3480 165 4050
rect 185 3480 200 4050
rect 150 3465 200 3480
rect 250 4050 300 4065
rect 250 3480 265 4050
rect 285 3480 300 4050
rect 250 3465 300 3480
rect 350 4050 400 4065
rect 350 3480 365 4050
rect 385 3480 400 4050
rect 350 3465 400 3480
rect 450 4050 500 4065
rect 450 3480 465 4050
rect 485 3480 500 4050
rect 450 3465 500 3480
rect 550 4050 600 4065
rect 550 3480 565 4050
rect 585 3480 600 4050
rect 550 3465 600 3480
rect -450 3275 -400 3290
rect -450 2105 -435 3275
rect -415 2105 -400 3275
rect -450 2090 -400 2105
rect -350 3275 -300 3290
rect -350 2105 -335 3275
rect -315 2105 -300 3275
rect -350 2090 -300 2105
rect -250 3275 -200 3290
rect -250 2105 -235 3275
rect -215 2105 -200 3275
rect -250 2090 -200 2105
rect -150 3275 -100 3290
rect -150 2105 -135 3275
rect -115 2105 -100 3275
rect -150 2090 -100 2105
rect -50 3275 0 3290
rect -50 2105 -35 3275
rect -15 2105 0 3275
rect -50 2090 0 2105
rect 50 3275 100 3290
rect 50 2105 65 3275
rect 85 2105 100 3275
rect 50 2090 100 2105
rect 150 3275 200 3290
rect 150 2105 165 3275
rect 185 2105 200 3275
rect 150 2090 200 2105
rect 250 3275 300 3290
rect 250 2105 265 3275
rect 285 2105 300 3275
rect 250 2090 300 2105
rect 350 3275 400 3290
rect 350 2105 365 3275
rect 385 2105 400 3275
rect 350 2090 400 2105
rect 450 3275 500 3290
rect 450 2105 465 3275
rect 485 2105 500 3275
rect 450 2090 500 2105
rect 550 3275 600 3290
rect 550 2105 565 3275
rect 585 2105 600 3275
rect 550 2090 600 2105
rect -450 1825 -400 1840
rect -450 1255 -435 1825
rect -415 1255 -400 1825
rect -450 1240 -400 1255
rect -350 1825 -300 1840
rect -350 1255 -335 1825
rect -315 1255 -300 1825
rect -350 1240 -300 1255
rect -250 1825 -200 1840
rect -250 1255 -235 1825
rect -215 1255 -200 1825
rect -250 1240 -200 1255
rect -150 1825 -100 1840
rect -150 1255 -135 1825
rect -115 1255 -100 1825
rect -150 1240 -100 1255
rect -50 1825 0 1840
rect -50 1255 -35 1825
rect -15 1255 0 1825
rect -50 1240 0 1255
rect 50 1825 100 1840
rect 50 1255 65 1825
rect 85 1255 100 1825
rect 50 1240 100 1255
rect 150 1825 200 1840
rect 150 1255 165 1825
rect 185 1255 200 1825
rect 150 1240 200 1255
rect 250 1825 300 1840
rect 250 1255 265 1825
rect 285 1255 300 1825
rect 250 1240 300 1255
rect 350 1825 400 1840
rect 350 1255 365 1825
rect 385 1255 400 1825
rect 350 1240 400 1255
rect 450 1825 500 1840
rect 450 1255 465 1825
rect 485 1255 500 1825
rect 450 1240 500 1255
rect 550 1825 600 1840
rect 550 1255 565 1825
rect 585 1255 600 1825
rect 550 1240 600 1255
<< ndiffc >>
rect -435 450 -415 1020
rect -335 450 -315 1020
rect -235 450 -215 1020
rect -135 450 -115 1020
rect -35 450 -15 1020
rect 65 450 85 1020
rect 165 450 185 1020
rect 265 450 285 1020
rect 365 450 385 1020
rect 465 450 485 1020
rect 565 450 585 1020
<< pdiffc >>
rect -435 3480 -415 4050
rect -335 3480 -315 4050
rect -235 3480 -215 4050
rect -135 3480 -115 4050
rect -35 3480 -15 4050
rect 65 3480 85 4050
rect 165 3480 185 4050
rect 265 3480 285 4050
rect 365 3480 385 4050
rect 465 3480 485 4050
rect 565 3480 585 4050
rect -435 2105 -415 3275
rect -335 2105 -315 3275
rect -235 2105 -215 3275
rect -135 2105 -115 3275
rect -35 2105 -15 3275
rect 65 2105 85 3275
rect 165 2105 185 3275
rect 265 2105 285 3275
rect 365 2105 385 3275
rect 465 2105 485 3275
rect 565 2105 585 3275
rect -435 1255 -415 1825
rect -335 1255 -315 1825
rect -235 1255 -215 1825
rect -135 1255 -115 1825
rect -35 1255 -15 1825
rect 65 1255 85 1825
rect 165 1255 185 1825
rect 265 1255 285 1825
rect 365 1255 385 1825
rect 465 1255 485 1825
rect 565 1255 585 1825
<< psubdiff >>
rect -500 1020 -450 1035
rect -500 450 -485 1020
rect -465 450 -450 1020
rect -500 435 -450 450
rect 600 1020 650 1035
rect 600 450 615 1020
rect 635 450 650 1020
rect 600 435 650 450
<< nsubdiff >>
rect -500 4050 -450 4065
rect -500 3480 -485 4050
rect -465 3480 -450 4050
rect -500 3465 -450 3480
rect 600 4050 650 4065
rect 600 3480 615 4050
rect 635 3480 650 4050
rect 600 3465 650 3480
rect -500 3275 -450 3290
rect -500 2105 -485 3275
rect -465 2105 -450 3275
rect -500 2090 -450 2105
rect 600 3275 650 3290
rect 600 2105 615 3275
rect 635 2105 650 3275
rect 600 2090 650 2105
rect -500 1825 -450 1840
rect -500 1255 -485 1825
rect -465 1255 -450 1825
rect -500 1240 -450 1255
rect 600 1825 650 1840
rect 600 1255 615 1825
rect 635 1255 650 1825
rect 600 1240 650 1255
<< psubdiffcont >>
rect -485 450 -465 1020
rect 615 450 635 1020
<< nsubdiffcont >>
rect -485 3480 -465 4050
rect 615 3480 635 4050
rect -485 2105 -465 3275
rect 615 2105 635 3275
rect -485 1255 -465 1825
rect 615 1255 635 1825
<< poly >>
rect -500 4150 450 4200
rect -450 4110 -350 4125
rect -450 4090 -435 4110
rect -415 4090 -350 4110
rect -450 4075 -350 4090
rect -400 4065 -350 4075
rect -300 4065 -250 4150
rect -200 4065 -150 4150
rect -100 4065 -50 4150
rect 0 4065 50 4150
rect 100 4065 150 4150
rect 200 4065 250 4150
rect 300 4065 350 4150
rect 400 4065 450 4150
rect 500 4110 600 4125
rect 500 4090 565 4110
rect 585 4090 600 4110
rect 500 4075 600 4090
rect 500 4065 550 4075
rect -400 3450 -350 3465
rect -300 3450 -250 3465
rect -200 3450 -150 3465
rect -100 3450 -50 3465
rect 0 3450 50 3465
rect 100 3450 150 3465
rect 200 3450 250 3465
rect 300 3450 350 3465
rect 400 3450 450 3465
rect 500 3450 550 3465
rect -500 3375 450 3425
rect -450 3335 -350 3350
rect -450 3315 -435 3335
rect -415 3315 -350 3335
rect -450 3300 -350 3315
rect -400 3290 -350 3300
rect -300 3290 -250 3375
rect -200 3290 -150 3375
rect -100 3290 -50 3305
rect 0 3290 50 3305
rect 100 3290 150 3305
rect 200 3290 250 3305
rect 300 3290 350 3375
rect 400 3290 450 3375
rect 500 3335 600 3350
rect 500 3315 565 3335
rect 585 3315 600 3335
rect 500 3300 600 3315
rect 500 3290 550 3300
rect -400 2075 -350 2090
rect -300 2075 -250 2090
rect -200 2075 -150 2090
rect -100 2050 -50 2090
rect 0 2050 50 2090
rect 100 2050 150 2090
rect 200 2050 250 2090
rect 300 2075 350 2090
rect 400 2075 450 2090
rect 500 2075 550 2090
rect -500 2000 250 2050
rect -500 1925 450 1975
rect -450 1885 -350 1900
rect -450 1865 -435 1885
rect -415 1865 -350 1885
rect -450 1850 -350 1865
rect -400 1840 -350 1850
rect -300 1840 -250 1925
rect -200 1840 -150 1855
rect -100 1840 -50 1855
rect 0 1840 50 1925
rect 100 1840 150 1925
rect 200 1840 250 1855
rect 300 1840 350 1855
rect 400 1840 450 1925
rect 500 1885 600 1900
rect 500 1865 565 1885
rect 585 1865 600 1885
rect 500 1850 600 1865
rect 500 1840 550 1850
rect -400 1225 -350 1240
rect -300 1225 -250 1240
rect -200 1200 -150 1240
rect -100 1200 -50 1240
rect 0 1225 50 1240
rect 100 1225 150 1240
rect 200 1200 250 1240
rect 300 1200 350 1240
rect 400 1225 450 1240
rect 500 1225 550 1240
rect -200 1185 350 1200
rect -200 1165 65 1185
rect 85 1165 350 1185
rect -200 1150 350 1165
rect -500 1075 450 1125
rect -400 1035 -350 1050
rect -300 1035 -250 1075
rect -200 1035 -150 1050
rect -100 1035 -50 1050
rect 0 1035 50 1075
rect 100 1035 150 1075
rect 200 1035 250 1050
rect 300 1035 350 1050
rect 400 1035 450 1075
rect 500 1035 550 1050
rect -400 425 -350 435
rect -450 410 -350 425
rect -300 420 -250 435
rect -450 390 -435 410
rect -415 390 -350 410
rect -450 375 -350 390
rect -200 350 -150 435
rect -100 350 -50 435
rect 0 420 50 435
rect 100 420 150 435
rect 200 350 250 435
rect 300 350 350 435
rect 400 420 450 435
rect 500 425 550 435
rect 500 410 600 425
rect 500 390 565 410
rect 585 390 600 410
rect 500 375 600 390
rect -500 300 350 350
<< polycont >>
rect -435 4090 -415 4110
rect 565 4090 585 4110
rect -435 3315 -415 3335
rect 565 3315 585 3335
rect -435 1865 -415 1885
rect 565 1865 585 1885
rect 65 1165 85 1185
rect -435 390 -415 410
rect 565 390 585 410
<< locali >>
rect -445 4110 -405 4120
rect -445 4090 -435 4110
rect -415 4090 -405 4110
rect -445 4060 -405 4090
rect 555 4110 595 4120
rect 555 4090 565 4110
rect 585 4090 595 4110
rect 555 4060 595 4090
rect -495 4050 -405 4060
rect -495 3480 -485 4050
rect -465 3480 -435 4050
rect -415 3480 -405 4050
rect -495 3470 -405 3480
rect -345 4050 -305 4060
rect -345 3480 -335 4050
rect -315 3480 -305 4050
rect -345 3470 -305 3480
rect -245 4050 -205 4060
rect -245 3480 -235 4050
rect -215 3480 -205 4050
rect -245 3470 -205 3480
rect -145 4050 -105 4060
rect -145 3480 -135 4050
rect -115 3480 -105 4050
rect -145 3445 -105 3480
rect -45 4050 -5 4060
rect -45 3480 -35 4050
rect -15 3480 -5 4050
rect -45 3470 -5 3480
rect 55 4050 95 4060
rect 55 3480 65 4050
rect 85 3480 95 4050
rect 55 3470 95 3480
rect 155 4050 195 4060
rect 155 3480 165 4050
rect 185 3480 195 4050
rect 155 3470 195 3480
rect 255 4050 295 4060
rect 255 3480 265 4050
rect 285 3480 295 4050
rect 255 3445 295 3480
rect 355 4050 395 4060
rect 355 3480 365 4050
rect 385 3480 395 4050
rect 355 3470 395 3480
rect 455 4050 495 4060
rect 455 3480 465 4050
rect 485 3480 495 4050
rect 455 3470 495 3480
rect 555 4050 645 4060
rect 555 3480 565 4050
rect 585 3480 615 4050
rect 635 3480 645 4050
rect 555 3470 645 3480
rect -145 3405 295 3445
rect -445 3335 -405 3345
rect -445 3315 -435 3335
rect -415 3315 -405 3335
rect -445 3285 -405 3315
rect -495 3275 -405 3285
rect -495 2105 -485 3275
rect -465 2105 -435 3275
rect -415 2105 -405 3275
rect -495 2095 -405 2105
rect -345 3275 -305 3285
rect -345 2105 -335 3275
rect -315 2105 -305 3275
rect -345 2095 -305 2105
rect -245 3275 -205 3285
rect -245 2105 -235 3275
rect -215 2105 -205 3275
rect -245 2095 -205 2105
rect -145 3275 -105 3405
rect -145 2105 -135 3275
rect -115 2105 -105 3275
rect -145 2095 -105 2105
rect -45 3275 -5 3285
rect -45 2105 -35 3275
rect -15 2105 -5 3275
rect -45 2095 -5 2105
rect 55 3275 95 3285
rect 55 2105 65 3275
rect 85 2105 95 3275
rect 55 2095 95 2105
rect 155 3275 195 3285
rect 155 2105 165 3275
rect 185 2105 195 3275
rect 155 2095 195 2105
rect 255 3275 295 3405
rect 555 3335 595 3345
rect 555 3315 565 3335
rect 585 3315 595 3335
rect 555 3285 595 3315
rect 255 2105 265 3275
rect 285 2105 295 3275
rect 255 2095 295 2105
rect 355 3275 395 3285
rect 355 2105 365 3275
rect 385 2105 395 3275
rect 355 2095 395 2105
rect 455 3275 495 3285
rect 455 2105 465 3275
rect 485 2105 495 3275
rect 455 2095 495 2105
rect 555 3275 645 3285
rect 555 2105 565 3275
rect 585 2105 615 3275
rect 635 2105 645 3275
rect 555 2095 645 2105
rect -445 1885 -405 1895
rect -445 1865 -435 1885
rect -415 1865 -405 1885
rect -445 1835 -405 1865
rect -495 1825 -405 1835
rect -495 1255 -485 1825
rect -465 1255 -435 1825
rect -415 1255 -405 1825
rect -495 1245 -405 1255
rect -345 1855 495 1895
rect -345 1825 -305 1855
rect -345 1255 -335 1825
rect -315 1255 -305 1825
rect -495 1020 -405 1030
rect -495 450 -485 1020
rect -465 450 -435 1020
rect -415 450 -405 1020
rect -495 440 -405 450
rect -445 410 -405 440
rect -445 390 -435 410
rect -415 390 -405 410
rect -445 380 -405 390
rect -345 1020 -305 1255
rect -245 1825 -205 1835
rect -245 1255 -235 1825
rect -215 1255 -205 1825
rect -245 1245 -205 1255
rect -145 1825 -105 1835
rect -145 1255 -135 1825
rect -115 1255 -105 1825
rect -145 1245 -105 1255
rect -45 1825 -5 1835
rect -45 1255 -35 1825
rect -15 1255 -5 1825
rect -45 1245 -5 1255
rect 55 1825 95 1835
rect 55 1255 65 1825
rect 85 1255 95 1825
rect 55 1185 95 1255
rect 155 1825 195 1835
rect 155 1255 165 1825
rect 185 1255 195 1825
rect 155 1245 195 1255
rect 255 1825 295 1835
rect 255 1255 265 1825
rect 285 1255 295 1825
rect 255 1245 295 1255
rect 355 1825 395 1835
rect 355 1255 365 1825
rect 385 1255 395 1825
rect 355 1245 395 1255
rect 455 1825 495 1855
rect 455 1255 465 1825
rect 485 1255 495 1825
rect 55 1165 65 1185
rect 85 1165 95 1185
rect -345 450 -335 1020
rect -315 450 -305 1020
rect -345 360 -305 450
rect -245 1020 -205 1030
rect -245 450 -235 1020
rect -215 450 -205 1020
rect -245 420 -205 450
rect -145 1020 -105 1030
rect -145 450 -135 1020
rect -115 450 -105 1020
rect -145 440 -105 450
rect -45 1020 -5 1030
rect -45 450 -35 1020
rect -15 450 -5 1020
rect -45 440 -5 450
rect 55 1020 95 1165
rect 455 1160 495 1255
rect 555 1885 595 1895
rect 555 1865 565 1885
rect 585 1865 595 1885
rect 555 1835 595 1865
rect 555 1825 645 1835
rect 555 1255 565 1825
rect 585 1255 615 1825
rect 635 1255 645 1825
rect 555 1245 645 1255
rect 455 1120 650 1160
rect 55 450 65 1020
rect 85 450 95 1020
rect 55 440 95 450
rect 155 1020 195 1030
rect 155 450 165 1020
rect 185 450 195 1020
rect 155 440 195 450
rect 255 1020 295 1030
rect 255 450 265 1020
rect 285 450 295 1020
rect 255 440 295 450
rect 355 1020 395 1030
rect 355 450 365 1020
rect 385 450 395 1020
rect 355 420 395 450
rect -245 380 395 420
rect 455 1020 495 1120
rect 455 450 465 1020
rect 485 450 495 1020
rect 455 360 495 450
rect 555 1020 645 1030
rect 555 450 565 1020
rect 585 450 615 1020
rect 635 450 645 1020
rect 555 440 645 450
rect 555 410 595 440
rect 555 390 565 410
rect 585 390 595 410
rect 555 380 595 390
rect -345 320 495 360
<< viali >>
rect -485 3480 -465 4050
rect -435 3480 -415 4050
rect -335 3480 -315 4050
rect 65 3480 85 4050
rect 465 3480 485 4050
rect 565 3480 585 4050
rect 615 3480 635 4050
rect -485 2105 -465 3275
rect -435 2105 -415 3275
rect -335 2105 -315 3275
rect 65 2105 85 3275
rect 465 2105 485 3275
rect 565 2105 585 3275
rect 615 2105 635 3275
rect -485 1255 -465 1825
rect -435 1255 -415 1825
rect -485 450 -465 1020
rect -435 450 -415 1020
rect -135 1255 -115 1825
rect 265 1255 285 1825
rect -235 450 -215 1020
rect -135 450 -115 1020
rect -35 450 -15 1020
rect 565 1255 585 1825
rect 615 1255 635 1825
rect 165 450 185 1020
rect 265 450 285 1020
rect 365 450 385 1020
rect 565 450 585 1020
rect 615 450 635 1020
<< metal1 >>
rect -500 4100 650 4250
rect -495 4050 -405 4100
rect -495 3480 -485 4050
rect -465 3480 -435 4050
rect -415 3480 -405 4050
rect -495 3275 -405 3480
rect -345 4050 -305 4100
rect -345 3480 -335 4050
rect -315 3480 -305 4050
rect -345 3470 -305 3480
rect -495 2105 -485 3275
rect -465 2105 -435 3275
rect -415 2105 -405 3275
rect -495 1825 -405 2105
rect -495 1255 -485 1825
rect -465 1255 -435 1825
rect -415 1255 -405 1825
rect -495 1245 -405 1255
rect -345 3275 -305 3285
rect -345 2105 -335 3275
rect -315 2105 -305 3275
rect -345 1160 -305 2105
rect -145 1825 -105 4100
rect 55 4050 95 4100
rect 55 3480 65 4050
rect 85 3480 95 4050
rect 55 3470 95 3480
rect 55 3275 95 3285
rect 55 2105 65 3275
rect 85 2105 95 3275
rect 55 2020 95 2105
rect -145 1255 -135 1825
rect -115 1255 -105 1825
rect -145 1245 -105 1255
rect -45 1970 195 2020
rect -345 1120 -205 1160
rect -495 1020 -405 1030
rect -495 450 -485 1020
rect -465 450 -435 1020
rect -415 450 -405 1020
rect -495 400 -405 450
rect -245 1020 -205 1120
rect -245 450 -235 1020
rect -215 450 -205 1020
rect -245 440 -205 450
rect -145 1020 -105 1030
rect -145 450 -135 1020
rect -115 450 -105 1020
rect -145 400 -105 450
rect -45 1020 -5 1970
rect -45 450 -35 1020
rect -15 450 -5 1020
rect -45 440 -5 450
rect 155 1020 195 1970
rect 255 1825 295 4100
rect 455 4050 495 4100
rect 455 3480 465 4050
rect 485 3480 495 4050
rect 455 3470 495 3480
rect 555 4050 645 4100
rect 555 3480 565 4050
rect 585 3480 615 4050
rect 635 3480 645 4050
rect 255 1255 265 1825
rect 285 1255 295 1825
rect 255 1245 295 1255
rect 455 3275 495 3285
rect 455 2105 465 3275
rect 485 2105 495 3275
rect 455 1160 495 2105
rect 555 3275 645 3480
rect 555 2105 565 3275
rect 585 2105 615 3275
rect 635 2105 645 3275
rect 555 1825 645 2105
rect 555 1255 565 1825
rect 585 1255 615 1825
rect 635 1255 645 1825
rect 555 1245 645 1255
rect 355 1120 495 1160
rect 155 450 165 1020
rect 185 450 195 1020
rect 155 440 195 450
rect 255 1020 295 1030
rect 255 450 265 1020
rect 285 450 295 1020
rect 255 400 295 450
rect 355 1020 395 1120
rect 355 450 365 1020
rect 385 450 395 1020
rect 355 440 395 450
rect 555 1020 645 1030
rect 555 450 565 1020
rect 585 450 615 1020
rect 635 450 645 1020
rect 555 400 645 450
rect -500 250 650 400
<< labels >>
rlabel metal1 -500 4170 -500 4170 3 VDD
rlabel poly -500 4175 -500 4175 7 Vbp
rlabel poly -500 3400 -500 3400 7 V2
rlabel pdiff -225 3465 -225 3465 5 net7
rlabel locali -125 4060 -125 4060 1 net8
rlabel poly -500 2025 -500 2025 7 V1
rlabel locali 375 3470 375 3470 5 net11
rlabel pdiff 175 2090 175 2090 5 net14
rlabel pdiff -25 2090 -25 2090 5 net13
rlabel pdiff -225 2090 -225 2090 5 net15
rlabel pdiff 375 2090 375 2090 5 net16
rlabel pdiff 375 1240 375 1240 5 net6
rlabel metal1 -500 285 -500 285 3 GND
rlabel poly -500 1950 -500 1950 7 Vcp
rlabel poly -500 1100 -500 1100 7 Vcn
rlabel poly -500 325 -500 325 7 Vbn
<< end >>
