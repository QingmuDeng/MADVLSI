magic
tech sky130A
timestamp 1615322015
<< error_p >>
rect -357 1160 -350 1200
rect -340 1143 -333 1217
rect 493 1143 500 1217
rect 510 1160 517 1200
<< nmos >>
rect -400 3465 -350 4065
rect -300 3465 -250 4065
rect -200 3465 -150 4065
rect -100 3465 -50 4065
rect 0 3465 50 4065
rect 100 3465 150 4065
rect 200 3465 250 4065
rect 300 3465 350 4065
rect 400 3465 450 4065
rect 500 3465 550 4065
rect -400 2065 -350 3265
rect -300 2065 -250 3265
rect -200 2065 -150 3265
rect -100 2065 -50 3265
rect 0 2065 50 3265
rect 100 2065 150 3265
rect 200 2065 250 3265
rect 300 2065 350 3265
rect 400 2065 450 3265
rect 500 2065 550 3265
rect -395 1215 -345 1815
rect -295 1215 -245 1815
rect -195 1215 -145 1815
rect -95 1215 -45 1815
rect 5 1215 55 1815
rect 105 1215 155 1815
rect 205 1215 255 1815
rect 305 1215 355 1815
rect 405 1215 455 1815
rect 505 1215 555 1815
rect -395 315 -345 915
rect -295 315 -245 915
rect -195 315 -145 915
rect -95 315 -45 915
rect 5 315 55 915
rect 105 315 155 915
rect 205 315 255 915
rect 305 315 355 915
rect 405 315 455 915
rect 505 315 555 915
<< ndiff >>
rect -450 4050 -400 4065
rect -450 3480 -435 4050
rect -415 3480 -400 4050
rect -450 3465 -400 3480
rect -350 4050 -300 4065
rect -350 3480 -335 4050
rect -315 3480 -300 4050
rect -350 3465 -300 3480
rect -250 4050 -200 4065
rect -250 3480 -235 4050
rect -215 3480 -200 4050
rect -250 3465 -200 3480
rect -150 4050 -100 4065
rect -150 3480 -135 4050
rect -115 3480 -100 4050
rect -150 3465 -100 3480
rect -50 4050 0 4065
rect -50 3480 -35 4050
rect -15 3480 0 4050
rect -50 3465 0 3480
rect 50 4050 100 4065
rect 50 3480 65 4050
rect 85 3480 100 4050
rect 50 3465 100 3480
rect 150 4050 200 4065
rect 150 3480 165 4050
rect 185 3480 200 4050
rect 150 3465 200 3480
rect 250 4050 300 4065
rect 250 3480 265 4050
rect 285 3480 300 4050
rect 250 3465 300 3480
rect 350 4050 400 4065
rect 350 3480 365 4050
rect 385 3480 400 4050
rect 350 3465 400 3480
rect 450 4050 500 4065
rect 450 3480 465 4050
rect 485 3480 500 4050
rect 450 3465 500 3480
rect 550 4050 600 4065
rect 550 3480 565 4050
rect 585 3480 600 4050
rect 550 3465 600 3480
rect -450 3250 -400 3265
rect -450 2080 -435 3250
rect -415 2080 -400 3250
rect -450 2065 -400 2080
rect -350 3250 -300 3265
rect -350 2080 -335 3250
rect -315 2080 -300 3250
rect -350 2065 -300 2080
rect -250 3250 -200 3265
rect -250 2080 -235 3250
rect -215 2080 -200 3250
rect -250 2065 -200 2080
rect -150 3250 -100 3265
rect -150 2080 -135 3250
rect -115 2080 -100 3250
rect -150 2065 -100 2080
rect -50 3250 0 3265
rect -50 2080 -35 3250
rect -15 2080 0 3250
rect -50 2065 0 2080
rect 50 3250 100 3265
rect 50 2080 65 3250
rect 85 2080 100 3250
rect 50 2065 100 2080
rect 150 3250 200 3265
rect 150 2080 165 3250
rect 185 2080 200 3250
rect 150 2065 200 2080
rect 250 3250 300 3265
rect 250 2080 265 3250
rect 285 2080 300 3250
rect 250 2065 300 2080
rect 350 3250 400 3265
rect 350 2080 365 3250
rect 385 2080 400 3250
rect 350 2065 400 2080
rect 450 3250 500 3265
rect 450 2080 465 3250
rect 485 2080 500 3250
rect 450 2065 500 2080
rect 550 3250 600 3265
rect 550 2080 565 3250
rect 585 2080 600 3250
rect 550 2065 600 2080
rect -445 1800 -395 1815
rect -445 1230 -430 1800
rect -410 1230 -395 1800
rect -445 1215 -395 1230
rect -345 1800 -295 1815
rect -345 1230 -330 1800
rect -310 1230 -295 1800
rect -345 1215 -295 1230
rect -245 1800 -195 1815
rect -245 1230 -230 1800
rect -210 1230 -195 1800
rect -245 1215 -195 1230
rect -145 1800 -95 1815
rect -145 1230 -130 1800
rect -110 1230 -95 1800
rect -145 1215 -95 1230
rect -45 1800 5 1815
rect -45 1230 -30 1800
rect -10 1230 5 1800
rect -45 1215 5 1230
rect 55 1800 105 1815
rect 55 1230 70 1800
rect 90 1230 105 1800
rect 55 1215 105 1230
rect 155 1800 205 1815
rect 155 1230 170 1800
rect 190 1230 205 1800
rect 155 1215 205 1230
rect 255 1800 305 1815
rect 255 1230 270 1800
rect 290 1230 305 1800
rect 255 1215 305 1230
rect 355 1800 405 1815
rect 355 1230 370 1800
rect 390 1230 405 1800
rect 355 1215 405 1230
rect 455 1800 505 1815
rect 455 1230 470 1800
rect 490 1230 505 1800
rect 455 1215 505 1230
rect 555 1800 605 1815
rect 555 1230 570 1800
rect 590 1230 605 1800
rect 555 1215 605 1230
rect -445 900 -395 915
rect -445 330 -430 900
rect -410 330 -395 900
rect -445 315 -395 330
rect -345 900 -295 915
rect -345 330 -330 900
rect -310 330 -295 900
rect -345 315 -295 330
rect -245 900 -195 915
rect -245 330 -230 900
rect -210 330 -195 900
rect -245 315 -195 330
rect -145 900 -95 915
rect -145 330 -130 900
rect -110 330 -95 900
rect -145 315 -95 330
rect -45 900 5 915
rect -45 330 -30 900
rect -10 330 5 900
rect -45 315 5 330
rect 55 900 105 915
rect 55 330 70 900
rect 90 330 105 900
rect 55 315 105 330
rect 155 900 205 915
rect 155 330 170 900
rect 190 330 205 900
rect 155 315 205 330
rect 255 900 305 915
rect 255 330 270 900
rect 290 330 305 900
rect 255 315 305 330
rect 355 900 405 915
rect 355 330 370 900
rect 390 330 405 900
rect 355 315 405 330
rect 455 900 505 915
rect 455 330 470 900
rect 490 330 505 900
rect 455 315 505 330
rect 555 900 605 915
rect 555 330 570 900
rect 590 330 605 900
rect 555 315 605 330
<< ndiffc >>
rect -435 3480 -415 4050
rect -335 3480 -315 4050
rect -235 3480 -215 4050
rect -135 3480 -115 4050
rect -35 3480 -15 4050
rect 65 3480 85 4050
rect 165 3480 185 4050
rect 265 3480 285 4050
rect 365 3480 385 4050
rect 465 3480 485 4050
rect 565 3480 585 4050
rect -435 2080 -415 3250
rect -335 2080 -315 3250
rect -235 2080 -215 3250
rect -135 2080 -115 3250
rect -35 2080 -15 3250
rect 65 2080 85 3250
rect 165 2080 185 3250
rect 265 2080 285 3250
rect 365 2080 385 3250
rect 465 2080 485 3250
rect 565 2080 585 3250
rect -430 1230 -410 1800
rect -330 1230 -310 1800
rect -230 1230 -210 1800
rect -130 1230 -110 1800
rect -30 1230 -10 1800
rect 70 1230 90 1800
rect 170 1230 190 1800
rect 270 1230 290 1800
rect 370 1230 390 1800
rect 470 1230 490 1800
rect 570 1230 590 1800
rect -430 330 -410 900
rect -330 330 -310 900
rect -230 330 -210 900
rect -130 330 -110 900
rect -30 330 -10 900
rect 70 330 90 900
rect 170 330 190 900
rect 270 330 290 900
rect 370 330 390 900
rect 470 330 490 900
rect 570 330 590 900
<< psubdiff >>
rect -500 4050 -450 4065
rect -500 3480 -485 4050
rect -465 3480 -450 4050
rect -500 3465 -450 3480
rect 600 4050 650 4065
rect 600 3480 615 4050
rect 635 3480 650 4050
rect 600 3465 650 3480
rect -500 3250 -450 3265
rect -500 2080 -485 3250
rect -465 2080 -450 3250
rect -500 2065 -450 2080
rect 600 3250 650 3265
rect 600 2080 615 3250
rect 635 2080 650 3250
rect 600 2065 650 2080
rect -495 1800 -445 1815
rect -495 1230 -480 1800
rect -460 1230 -445 1800
rect -495 1215 -445 1230
rect 605 1800 655 1815
rect 605 1230 620 1800
rect 640 1230 655 1800
rect 605 1215 655 1230
rect -495 900 -445 915
rect -495 330 -480 900
rect -460 330 -445 900
rect -495 315 -445 330
rect 605 900 655 915
rect 605 330 620 900
rect 640 330 655 900
rect 605 315 655 330
<< psubdiffcont >>
rect -485 3480 -465 4050
rect 615 3480 635 4050
rect -485 2080 -465 3250
rect 615 2080 635 3250
rect -480 1230 -460 1800
rect 620 1230 640 1800
rect -480 330 -460 900
rect 620 330 640 900
<< poly >>
rect -400 4110 -350 4125
rect -400 4090 -385 4110
rect -365 4090 -350 4110
rect -400 4065 -350 4090
rect -300 4110 -250 4125
rect -300 4090 -285 4110
rect -265 4090 -250 4110
rect -300 4065 -250 4090
rect -200 4110 -150 4125
rect -200 4090 -185 4110
rect -165 4090 -150 4110
rect -200 4065 -150 4090
rect -100 4110 -50 4125
rect -100 4090 -85 4110
rect -65 4090 -50 4110
rect -100 4065 -50 4090
rect 0 4110 50 4125
rect 0 4090 15 4110
rect 35 4090 50 4110
rect 0 4065 50 4090
rect 100 4110 150 4125
rect 100 4090 115 4110
rect 135 4090 150 4110
rect 100 4065 150 4090
rect 200 4110 250 4125
rect 200 4090 215 4110
rect 235 4090 250 4110
rect 200 4065 250 4090
rect 300 4110 350 4125
rect 300 4090 315 4110
rect 335 4090 350 4110
rect 300 4065 350 4090
rect 400 4110 450 4125
rect 400 4090 415 4110
rect 435 4090 450 4110
rect 400 4065 450 4090
rect 500 4110 550 4125
rect 500 4090 515 4110
rect 535 4090 550 4110
rect 500 4065 550 4090
rect -400 3450 -350 3465
rect -300 3450 -250 3465
rect -200 3450 -150 3465
rect -100 3450 -50 3465
rect 0 3450 50 3465
rect 100 3450 150 3465
rect 200 3450 250 3465
rect 300 3450 350 3465
rect 400 3450 450 3465
rect 500 3450 550 3465
rect -400 3310 -350 3325
rect -400 3290 -385 3310
rect -365 3290 -350 3310
rect -400 3265 -350 3290
rect -300 3310 450 3345
rect -300 3290 -285 3310
rect -265 3305 450 3310
rect -265 3290 -250 3305
rect -300 3265 -250 3290
rect -200 3265 -150 3305
rect -100 3265 -50 3280
rect 0 3265 50 3280
rect 100 3265 150 3280
rect 200 3265 250 3280
rect 300 3265 350 3305
rect 400 3265 450 3305
rect 500 3310 550 3325
rect 500 3290 515 3310
rect 535 3290 550 3310
rect 500 3265 550 3290
rect -400 2050 -350 2065
rect -300 2050 -250 2065
rect -200 2050 -150 2065
rect -100 2050 -50 2065
rect 0 2050 50 2065
rect 100 2050 150 2065
rect 200 2050 250 2065
rect 300 2050 350 2065
rect 400 2050 450 2065
rect 500 2050 550 2065
rect -100 2005 250 2050
rect -195 1855 355 1905
rect -395 1815 -345 1830
rect -295 1815 -245 1830
rect -195 1815 -145 1855
rect -95 1815 -45 1855
rect 5 1815 55 1830
rect 105 1815 155 1830
rect 205 1815 255 1855
rect 305 1815 355 1855
rect 405 1815 455 1830
rect 505 1815 555 1830
rect -395 1190 -345 1215
rect -395 1170 -380 1190
rect -360 1170 -345 1190
rect -395 1155 -345 1170
rect -295 1175 -245 1215
rect -195 1200 -145 1215
rect -95 1200 -45 1215
rect 5 1175 55 1215
rect 105 1175 155 1215
rect 205 1200 255 1215
rect 305 1200 355 1215
rect 405 1175 455 1215
rect 505 1190 555 1215
rect -295 1125 460 1175
rect 505 1170 520 1190
rect 540 1170 555 1190
rect 505 1155 555 1170
rect -195 955 355 1005
rect -395 915 -345 930
rect -295 915 -245 930
rect -195 915 -145 955
rect -95 915 -45 955
rect 5 915 55 930
rect 105 915 155 930
rect 205 915 255 955
rect 305 915 355 955
rect 405 915 455 930
rect 505 915 555 930
rect -395 290 -345 315
rect -395 270 -380 290
rect -360 270 -345 290
rect -395 255 -345 270
rect -295 275 -245 315
rect -195 300 -145 315
rect -95 300 -45 315
rect 5 275 55 315
rect 105 275 155 315
rect 205 300 255 315
rect 305 300 355 315
rect 405 275 455 315
rect -295 225 455 275
rect 505 290 555 315
rect 505 270 520 290
rect 540 270 555 290
rect 505 255 555 270
<< polycont >>
rect -385 4090 -365 4110
rect -285 4090 -265 4110
rect -185 4090 -165 4110
rect -85 4090 -65 4110
rect 15 4090 35 4110
rect 115 4090 135 4110
rect 215 4090 235 4110
rect 315 4090 335 4110
rect 415 4090 435 4110
rect 515 4090 535 4110
rect -385 3290 -365 3310
rect -285 3290 -265 3310
rect 515 3290 535 3310
rect -380 1170 -360 1190
rect 520 1170 540 1190
rect -380 270 -360 290
rect 520 270 540 290
<< locali >>
rect -395 4110 545 4120
rect -395 4090 -385 4110
rect -365 4090 -285 4110
rect -265 4090 -185 4110
rect -165 4090 -85 4110
rect -65 4090 15 4110
rect 35 4090 115 4110
rect 135 4090 215 4110
rect 235 4090 315 4110
rect 335 4090 415 4110
rect 435 4090 515 4110
rect 535 4090 545 4110
rect -395 4080 545 4090
rect -495 4050 -405 4060
rect -495 3480 -485 4050
rect -465 3480 -435 4050
rect -415 3480 -405 4050
rect -495 3470 -405 3480
rect -345 4050 -305 4060
rect -345 3480 -335 4050
rect -315 3480 -305 4050
rect -345 3470 -305 3480
rect -245 4050 -205 4060
rect -245 3480 -235 4050
rect -215 3480 -205 4050
rect -245 3470 -205 3480
rect -145 4050 -105 4060
rect -145 3480 -135 4050
rect -115 3480 -105 4050
rect -145 3445 -105 3480
rect -45 4050 -5 4060
rect -45 3480 -35 4050
rect -15 3480 -5 4050
rect -45 3470 -5 3480
rect 55 4050 95 4060
rect 55 3480 65 4050
rect 85 3480 95 4050
rect 55 3470 95 3480
rect 155 4050 195 4060
rect 155 3480 165 4050
rect 185 3480 195 4050
rect 155 3470 195 3480
rect 255 4050 295 4060
rect 255 3480 265 4050
rect 285 3480 295 4050
rect 255 3445 295 3480
rect 355 4050 395 4060
rect 355 3480 365 4050
rect 385 3480 395 4050
rect 355 3470 395 3480
rect 455 4050 495 4060
rect 455 3480 465 4050
rect 485 3480 495 4050
rect 455 3470 495 3480
rect 555 4050 645 4060
rect 555 3480 565 4050
rect 585 3480 615 4050
rect 635 3480 645 4050
rect 555 3470 645 3480
rect -145 3405 295 3445
rect -395 3310 -355 3320
rect -395 3290 -385 3310
rect -365 3290 -355 3310
rect -395 3280 -355 3290
rect -295 3310 -255 3320
rect -295 3290 -285 3310
rect -265 3290 -255 3310
rect -295 3280 -255 3290
rect -495 3250 -405 3260
rect -495 2080 -485 3250
rect -465 2080 -435 3250
rect -415 2080 -405 3250
rect -495 2070 -405 2080
rect -345 3250 -305 3260
rect -345 2080 -335 3250
rect -315 2080 -305 3250
rect -345 2070 -305 2080
rect -245 3250 -205 3260
rect -245 2080 -235 3250
rect -215 2080 -205 3250
rect -245 2070 -205 2080
rect -145 3250 -105 3405
rect -145 2080 -135 3250
rect -115 2080 -105 3250
rect -145 2070 -105 2080
rect -45 3250 -5 3260
rect -45 2080 -35 3250
rect -15 2080 -5 3250
rect -45 2070 -5 2080
rect 55 3250 95 3265
rect 55 2080 65 3250
rect 85 2080 95 3250
rect 55 1965 95 2080
rect 155 3250 195 3260
rect 155 2080 165 3250
rect 185 2080 195 3250
rect 155 2070 195 2080
rect 255 3250 295 3405
rect 505 3310 545 3320
rect 505 3290 515 3310
rect 535 3290 545 3310
rect 505 3280 545 3290
rect 255 2080 265 3250
rect 285 2080 295 3250
rect 255 2070 295 2080
rect 355 3250 395 3260
rect 355 2080 365 3250
rect 385 2080 395 3250
rect 355 2070 395 2080
rect 455 3250 495 3260
rect 455 2080 465 3250
rect 485 2080 495 3250
rect 455 2070 495 2080
rect 555 3250 645 3260
rect 555 2080 565 3250
rect 585 2080 615 3250
rect 635 2080 645 3250
rect 555 2070 645 2080
rect -490 1800 -400 1810
rect -490 1230 -480 1800
rect -460 1230 -430 1800
rect -410 1230 -400 1800
rect -490 1220 -400 1230
rect -340 1800 -300 1810
rect -340 1230 -330 1800
rect -310 1230 -300 1800
rect -340 1200 -300 1230
rect -240 1800 -200 1810
rect -240 1230 -230 1800
rect -210 1230 -200 1800
rect -240 1220 -200 1230
rect -140 1800 -100 1810
rect -140 1230 -130 1800
rect -110 1230 -100 1800
rect -140 1220 -100 1230
rect -40 1800 0 1810
rect -40 1230 -30 1800
rect -10 1230 0 1800
rect -40 1220 0 1230
rect 60 1800 100 1830
rect 60 1230 70 1800
rect 90 1230 100 1800
rect 60 1220 100 1230
rect 160 1800 200 1810
rect 160 1230 170 1800
rect 190 1230 200 1800
rect 160 1220 200 1230
rect 260 1800 300 1810
rect 260 1230 270 1800
rect 290 1230 300 1800
rect 260 1220 300 1230
rect 360 1800 400 1810
rect 360 1230 370 1800
rect 390 1230 400 1800
rect 360 1220 400 1230
rect 460 1800 500 1810
rect 460 1230 470 1800
rect 490 1230 500 1800
rect 460 1200 500 1230
rect 560 1800 650 1810
rect 560 1230 570 1800
rect 590 1230 620 1800
rect 640 1230 650 1800
rect 560 1220 650 1230
rect -390 1190 -350 1200
rect -390 1170 -380 1190
rect -360 1170 -350 1190
rect -390 1160 -350 1170
rect -340 1160 500 1200
rect 510 1190 550 1200
rect 510 1170 520 1190
rect 540 1170 550 1190
rect 510 1160 550 1170
rect -490 900 -400 910
rect -490 330 -480 900
rect -460 330 -430 900
rect -410 330 -400 900
rect -490 320 -400 330
rect -340 900 -300 1160
rect -340 330 -330 900
rect -310 330 -300 900
rect -340 320 -300 330
rect -240 900 -200 910
rect -240 330 -230 900
rect -210 330 -200 900
rect -240 320 -200 330
rect -140 900 -100 910
rect -140 330 -130 900
rect -110 330 -100 900
rect -140 320 -100 330
rect -40 900 0 910
rect -40 330 -30 900
rect -10 330 0 900
rect -40 320 0 330
rect 60 900 100 910
rect 60 330 70 900
rect 90 330 100 900
rect 60 320 100 330
rect 160 900 200 910
rect 160 330 170 900
rect 190 330 200 900
rect 160 320 200 330
rect 260 900 300 910
rect 260 330 270 900
rect 290 330 300 900
rect 260 320 300 330
rect 360 900 400 910
rect 360 330 370 900
rect 390 330 400 900
rect 360 320 400 330
rect 460 900 500 1160
rect 460 330 470 900
rect 490 330 500 900
rect 460 320 500 330
rect 560 900 650 910
rect 560 330 570 900
rect 590 330 620 900
rect 640 330 650 900
rect 560 320 650 330
rect -390 290 -350 300
rect -390 270 -380 290
rect -360 270 -350 290
rect -390 260 -350 270
rect 510 290 550 300
rect 510 270 520 290
rect 540 270 550 290
rect 510 260 550 270
<< end >>
