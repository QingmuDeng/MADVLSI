magic
tech sky130A
timestamp 1614097730
<< nwell >>
rect -145 500 20 915
<< nmos >>
rect -75 365 -60 465
<< pmos >>
rect -75 795 -60 895
<< ndiff >>
rect -125 450 -75 465
rect -125 380 -110 450
rect -90 380 -75 450
rect -125 365 -75 380
rect -60 450 -10 465
rect -60 380 -45 450
rect -25 380 -10 450
rect -60 365 -10 380
<< pdiff >>
rect -125 880 -75 895
rect -125 810 -110 880
rect -90 810 -75 880
rect -125 795 -75 810
rect -60 880 -10 895
rect -60 810 -45 880
rect -25 810 -10 880
rect -60 795 -10 810
<< ndiffc >>
rect -110 380 -90 450
rect -45 380 -25 450
<< pdiffc >>
rect -110 810 -90 880
rect -45 810 -25 880
<< psubdiff >>
rect -125 310 -75 325
rect -125 240 -110 310
rect -90 240 -75 310
rect -125 225 -75 240
<< nsubdiff >>
rect -50 715 0 730
rect -50 645 -35 715
rect -15 645 0 715
rect -50 630 0 645
<< psubdiffcont >>
rect -110 240 -90 310
<< nsubdiffcont >>
rect -35 645 -15 715
<< poly >>
rect -100 940 -60 950
rect -100 920 -90 940
rect -70 920 -60 940
rect -100 910 -60 920
rect -75 895 -60 910
rect -75 615 -60 795
rect -75 605 -35 615
rect -75 585 -65 605
rect -45 585 -35 605
rect -75 575 -35 585
rect -75 465 -60 575
rect -75 350 -60 365
<< polycont >>
rect -90 920 -70 940
rect -65 585 -45 605
<< locali >>
rect -100 940 -60 950
rect -100 930 -90 940
rect -145 920 -90 930
rect -70 920 -60 940
rect -145 910 -60 920
rect -120 880 -80 890
rect -120 810 -110 880
rect -90 810 -80 880
rect -120 800 -80 810
rect -55 880 -15 890
rect -55 810 -45 880
rect -25 820 -15 880
rect -25 810 5 820
rect -55 800 5 810
rect -35 765 -15 800
rect -120 745 -15 765
rect -120 460 -100 745
rect -45 715 -5 725
rect -45 645 -35 715
rect -15 645 -5 715
rect -45 635 -5 645
rect -75 605 5 615
rect -75 585 -65 605
rect -45 595 5 605
rect -45 585 -35 595
rect -75 575 -35 585
rect -120 450 -80 460
rect -120 380 -110 450
rect -90 380 -80 450
rect -120 370 -80 380
rect -55 450 -15 460
rect -55 380 -45 450
rect -25 380 -15 450
rect -55 370 -15 380
rect -120 310 -80 320
rect -120 240 -110 310
rect -90 240 -80 310
rect -120 230 -80 240
<< viali >>
rect -110 810 -90 880
rect -35 645 -15 715
rect -45 380 -25 450
rect -110 240 -90 310
<< metal1 >>
rect -145 880 5 895
rect -145 810 -110 880
rect -90 810 5 880
rect -145 715 5 810
rect -145 645 -35 715
rect -15 645 5 715
rect -145 520 5 645
rect -145 450 5 465
rect -145 380 -45 450
rect -25 380 5 450
rect -145 310 5 380
rect -145 240 -110 310
rect -90 240 5 310
rect -145 90 5 240
rect -145 -5 5 35
<< labels >>
rlabel locali -145 920 -145 920 7 D
port 1 w
rlabel metal1 -145 715 -145 715 7 VP
port 3 w
rlabel metal1 -145 265 -145 265 7 VN
port 4 w
rlabel metal1 -145 15 -145 15 7 CLK
port 2 w
rlabel locali 5 810 5 810 3 nD
port 5 e
<< end >>
