magic
tech sky130A
timestamp 1615758221
<< poly >>
rect 3215 3110 3385 3160
rect 3215 3010 3265 3110
rect 3215 2980 3225 3010
rect 3255 2980 3265 3010
rect 3215 2970 3265 2980
rect 3165 2335 3375 2385
rect 3165 1735 3215 2335
rect 3165 1705 3175 1735
rect 3205 1705 3215 1735
rect 3165 1695 3215 1705
rect 3165 1595 3215 1605
rect 3165 1565 3175 1595
rect 3205 1565 3215 1595
rect 3165 1010 3215 1565
rect 3165 960 3400 1010
rect 3215 925 3285 935
rect 3215 895 3225 925
rect 3255 895 3285 925
rect 3215 885 3285 895
rect 3215 75 3285 85
rect 3215 45 3225 75
rect 3255 45 3285 75
rect 3215 35 3285 45
rect 3215 -565 3265 -555
rect 3215 -595 3225 -565
rect 3255 -595 3265 -565
rect 3215 -690 3265 -595
rect 3215 -740 3285 -690
<< polycont >>
rect 3225 2980 3255 3010
rect 3175 1705 3205 1735
rect 3175 1565 3205 1595
rect 3225 895 3255 925
rect 3225 45 3255 75
rect 3225 -595 3255 -565
<< locali >>
rect 3215 3010 3265 3020
rect 3215 2980 3225 3010
rect 3255 2980 3265 3010
rect 3215 2970 3265 2980
rect 2735 1780 3215 1830
rect 2735 1710 3145 1760
rect 3095 1605 3145 1710
rect 3165 1735 3215 1780
rect 3165 1705 3175 1735
rect 3205 1705 3215 1735
rect 3165 1695 3215 1705
rect 3095 1595 3215 1605
rect 3095 1565 3175 1595
rect 3205 1565 3215 1595
rect 3095 1555 3215 1565
rect 3215 925 3265 935
rect 3215 895 3225 925
rect 3255 895 3265 925
rect 3215 885 3265 895
rect 3215 75 3265 85
rect 3215 45 3225 75
rect 3255 45 3265 75
rect 3215 35 3265 45
rect 3215 -565 3265 -555
rect 3215 -595 3225 -565
rect 3255 -595 3265 -565
rect 3215 -605 3265 -595
<< viali >>
rect 3225 2980 3255 3010
rect 3225 895 3255 925
rect 3225 45 3255 75
rect 3225 -595 3255 -565
<< metal1 >>
rect 2780 3060 3405 3210
rect 2780 1040 3100 3060
rect 3215 3010 3265 3020
rect 3215 2980 3225 3010
rect 3255 2980 3265 3010
rect 3215 1010 3265 2980
rect 2905 960 3265 1010
rect 2940 925 3265 935
rect 2940 895 3225 925
rect 3255 895 3265 925
rect 2940 885 3265 895
rect 2940 810 3265 860
rect 2940 730 3190 780
rect 2780 -640 3105 700
rect 3140 10 3190 730
rect 3215 75 3265 810
rect 3215 45 3225 75
rect 3255 45 3265 75
rect 3215 35 3265 45
rect 3140 -40 3265 10
rect 3215 -565 3265 -40
rect 3215 -595 3225 -565
rect 3255 -595 3265 -565
rect 3215 -605 3265 -595
rect 2780 -790 3440 -640
use cas_diff_lvs  cas_diff_lvs_0
timestamp 1615756184
transform 1 0 3785 0 1 -1040
box -520 250 670 4250
use bias_lvs  bias_lvs_0
timestamp 1615435668
transform 1 0 2424 0 1 -275
box -2415 285 580 2005
<< end >>
