* SPICE3 file created from /home/madvlsi/MADVLSI/mini3/layout/cas_diff_lvs.ext - technology: sky130A


* Top level circuit /home/madvlsi/MADVLSI/mini3/layout/cas_diff_lvs

X0 a_n700_880# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=6e+12p pd=2.6e+07u as=3.9e+13p ps=1.67e+08u w=6e+06u l=500000u
X1 net6 a_n400_2310# VDD VDD sky130_fd_pr__pfet_01v8 ad=3e+12p pd=1.3e+07u as=0p ps=0u w=6e+06u l=500000u
X2 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=500000u
X3 a_n700_4180# Vcn a_n700_880# GND sky130_fd_pr__nfet_01v8 ad=6e+12p pd=2.6e+07u as=6e+12p ps=2.6e+07u w=6e+06u l=500000u
X4 a_n400_2310# Vcn a_n100_880# GND sky130_fd_pr__nfet_01v8 ad=3e+12p pd=1.3e+07u as=6e+12p ps=2.6e+07u w=6e+06u l=500000u
X5 net8 V2 net15 VDD sky130_fd_pr__pfet_01v8 ad=1.8e+13p pd=7.6e+07u as=6e+12p ps=2.5e+07u w=1.2e+07u l=500000u
X6 net14 V1 a_n100_880# VDD sky130_fd_pr__pfet_01v8 ad=6e+12p pd=2.5e+07u as=6e+12p ps=2.5e+07u w=1.2e+07u l=500000u
X7 a_n700_880# Vcn a_n700_4180# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=500000u
X8 GND GND a_n700_880# GND sky130_fd_pr__nfet_01v8 ad=1.2e+13p pd=5.2e+07u as=0p ps=0u w=6e+06u l=500000u
X9 net7 Vbp VDD VDD sky130_fd_pr__pfet_01v8 ad=3e+12p pd=1.3e+07u as=0p ps=0u w=6e+06u l=500000u
X10 net8 Vbp a_300_6930# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3e+12p ps=1.3e+07u w=6e+06u l=500000u
X11 VDD VDD a_n700_880# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=500000u
X12 a_n100_880# Vbn GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=500000u
X13 a_n500_2490# Vcp a_n700_880# VDD sky130_fd_pr__pfet_01v8 ad=3e+12p pd=1.3e+07u as=0p ps=0u w=6e+06u l=500000u
X14 VDD a_n400_2310# a_300_2490# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3e+12p ps=1.3e+07u w=6e+06u l=500000u
X15 GND Vbn a_n100_880# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=500000u
X16 a_n700_4180# V2 net16 VDD sky130_fd_pr__pfet_01v8 ad=1.2e+13p pd=5e+07u as=6e+12p ps=2.5e+07u w=1.2e+07u l=500000u
X17 net13 V1 net8 VDD sky130_fd_pr__pfet_01v8 ad=6e+12p pd=2.5e+07u as=0p ps=0u w=1.2e+07u l=500000u
X18 net8 Vbp net7 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=500000u
X19 a_300_6930# Vbp VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=500000u
X20 a_n100_880# V1 net13 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.2e+07u l=500000u
X21 a_n700_880# GND GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=500000u
X22 VDD a_n400_2310# a_n500_2490# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=500000u
X23 a_300_2490# Vcp a_n400_2310# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3e+12p ps=1.3e+07u w=6e+06u l=500000u
X24 a_n700_4180# VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.2e+07u l=500000u
X25 net16 V2 net8 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.2e+07u l=500000u
X26 VDD Vbp net11 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3e+12p ps=1.3e+07u w=6e+06u l=500000u
X27 GND Vbn a_n700_4180# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=500000u
X28 a_n100_6930# Vbp net8 VDD sky130_fd_pr__pfet_01v8 ad=3e+12p pd=1.3e+07u as=0p ps=0u w=6e+06u l=500000u
X29 VDD VDD a_n700_4180# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.2e+07u l=500000u
X30 a_n700_4180# Vbn GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=500000u
X31 a_n700_880# Vcp net6 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=500000u
X32 VDD Vbp a_n100_6930# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=500000u
X33 a_n100_2490# a_n400_2310# VDD VDD sky130_fd_pr__pfet_01v8 ad=3e+12p pd=1.3e+07u as=0p ps=0u w=6e+06u l=500000u
X34 net15 V2 a_n700_4180# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.2e+07u l=500000u
X35 net8 V1 net14 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.2e+07u l=500000u
X36 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=500000u
X37 net11 Vbp net8 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=500000u
X38 a_n100_880# Vcn a_n400_2310# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=500000u
X39 a_n400_2310# Vcp a_n100_2490# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=6e+06u l=500000u
.end

