magic
tech sky130A
timestamp 1613924644
<< nwell >>
rect -85 195 255 645
<< nmos >>
rect 0 -5 15 95
rect 40 -5 55 95
rect 105 -5 120 95
rect 170 -5 185 95
rect 0 -280 15 -180
rect 40 -280 55 -180
rect 105 -280 120 -180
rect 170 -280 185 -180
<< pmos >>
rect 0 490 15 590
rect 65 490 80 590
rect 130 490 145 590
rect 170 490 185 590
rect 0 215 15 315
rect 65 215 80 315
rect 130 215 145 315
rect 170 215 185 315
<< ndiff >>
rect -50 80 0 95
rect -50 10 -35 80
rect -15 10 0 80
rect -50 -5 0 10
rect 15 -5 40 95
rect 55 80 105 95
rect 55 10 70 80
rect 90 10 105 80
rect 55 -5 105 10
rect 120 80 170 95
rect 120 10 135 80
rect 155 10 170 80
rect 120 -5 170 10
rect 185 80 235 95
rect 185 10 200 80
rect 220 10 235 80
rect 185 -5 235 10
rect -50 -195 0 -180
rect -50 -265 -35 -195
rect -15 -265 0 -195
rect -50 -280 0 -265
rect 15 -280 40 -180
rect 55 -195 105 -180
rect 55 -265 70 -195
rect 90 -265 105 -195
rect 55 -280 105 -265
rect 120 -195 170 -180
rect 120 -265 135 -195
rect 155 -265 170 -195
rect 120 -280 170 -265
rect 185 -195 235 -180
rect 185 -265 200 -195
rect 220 -265 235 -195
rect 185 -280 235 -265
<< pdiff >>
rect -50 575 0 590
rect -50 505 -35 575
rect -15 505 0 575
rect -50 490 0 505
rect 15 575 65 590
rect 15 505 30 575
rect 50 505 65 575
rect 15 490 65 505
rect 80 575 130 590
rect 80 505 95 575
rect 115 505 130 575
rect 80 490 130 505
rect 145 490 170 590
rect 185 575 235 590
rect 185 505 200 575
rect 220 505 235 575
rect 185 490 235 505
rect -50 300 0 315
rect -50 230 -35 300
rect -15 230 0 300
rect -50 215 0 230
rect 15 300 65 315
rect 15 230 30 300
rect 50 230 65 300
rect 15 215 65 230
rect 80 300 130 315
rect 80 230 95 300
rect 115 230 130 300
rect 80 215 130 230
rect 145 215 170 315
rect 185 300 235 315
rect 185 230 200 300
rect 220 230 235 300
rect 185 215 235 230
<< ndiffc >>
rect -35 10 -15 80
rect 70 10 90 80
rect 135 10 155 80
rect 200 10 220 80
rect -35 -265 -15 -195
rect 70 -265 90 -195
rect 135 -265 155 -195
rect 200 -265 220 -195
<< pdiffc >>
rect -35 505 -15 575
rect 30 505 50 575
rect 95 505 115 575
rect 200 505 220 575
rect -35 230 -15 300
rect 30 230 50 300
rect 95 230 115 300
rect 200 230 220 300
<< psubdiff >>
rect -65 -60 -15 -45
rect -65 -130 -50 -60
rect -30 -130 -15 -60
rect -65 -145 -15 -130
<< nsubdiff >>
rect -60 440 -10 455
rect -60 370 -45 440
rect -25 370 -10 440
rect -60 355 -10 370
<< psubdiffcont >>
rect -50 -130 -30 -60
<< nsubdiffcont >>
rect -45 370 -25 440
<< poly >>
rect 170 605 210 645
rect 0 590 15 605
rect 65 590 80 605
rect 130 590 145 605
rect 170 590 185 605
rect 0 315 15 490
rect 65 475 80 490
rect 65 435 105 475
rect 40 370 80 410
rect 65 315 80 370
rect 130 315 145 490
rect 170 475 185 490
rect 190 390 230 430
rect 210 340 230 390
rect 170 325 230 340
rect 170 315 185 325
rect 0 200 15 215
rect 65 200 80 215
rect 130 200 145 215
rect 170 200 185 215
rect 0 95 15 110
rect 40 95 55 110
rect 105 95 120 110
rect 170 95 185 110
rect 0 -180 15 -5
rect 40 -75 55 -5
rect 40 -115 80 -75
rect 40 -180 55 -165
rect 105 -180 120 -5
rect 170 -60 185 -5
rect 145 -100 185 -60
rect 170 -165 210 -125
rect 170 -180 185 -165
rect 0 -295 15 -280
rect 40 -295 55 -280
rect 105 -295 120 -280
rect 170 -295 185 -280
rect 40 -335 80 -295
<< locali >>
rect 170 625 210 645
rect 145 605 210 625
rect -45 575 -5 585
rect -45 505 -35 575
rect -15 505 -5 575
rect -45 495 -5 505
rect 20 575 60 585
rect 20 505 30 575
rect 50 505 60 575
rect 20 495 60 505
rect 85 575 125 585
rect 85 505 95 575
rect 115 505 125 575
rect 85 495 125 505
rect -55 440 -15 450
rect -55 370 -45 440
rect -25 370 -15 440
rect 20 410 40 495
rect 65 455 105 475
rect 65 435 120 455
rect 20 390 80 410
rect 40 370 80 390
rect -55 360 -15 370
rect 100 350 120 435
rect 40 330 120 350
rect 40 310 60 330
rect 145 310 165 605
rect 190 575 230 585
rect 190 505 200 575
rect 220 505 230 575
rect 190 495 230 505
rect 210 430 230 495
rect 190 390 230 430
rect -45 300 -5 310
rect -45 230 -35 300
rect -15 230 -5 300
rect -45 220 -5 230
rect 20 300 60 310
rect 20 230 30 300
rect 50 230 60 300
rect 20 220 60 230
rect 85 300 125 310
rect 85 230 95 300
rect 115 230 125 300
rect 145 300 230 310
rect 145 290 200 300
rect 85 220 125 230
rect 190 230 200 290
rect 220 230 230 300
rect 190 220 230 230
rect -45 80 -5 90
rect -45 10 -35 80
rect -15 10 -5 80
rect 60 80 100 90
rect 60 20 70 80
rect -45 0 -5 10
rect 15 10 70 20
rect 90 10 100 80
rect 15 0 100 10
rect 125 80 165 90
rect 125 10 135 80
rect 155 10 165 80
rect 125 0 165 10
rect 190 80 230 90
rect 190 10 200 80
rect 220 10 230 80
rect 190 0 230 10
rect 15 -20 35 0
rect 0 -40 35 -20
rect 145 -20 165 0
rect 145 -40 225 -20
rect -60 -60 -20 -50
rect -60 -130 -50 -60
rect -30 -130 -20 -60
rect -60 -140 -20 -130
rect 0 -145 20 -40
rect 40 -115 80 -75
rect 145 -80 185 -60
rect 0 -165 35 -145
rect -45 -195 -5 -185
rect -45 -265 -35 -195
rect -15 -265 -5 -195
rect -45 -275 -5 -265
rect 15 -295 35 -165
rect 60 -185 80 -115
rect 125 -100 185 -80
rect 125 -185 145 -100
rect 205 -125 225 -40
rect 170 -145 225 -125
rect 170 -165 210 -145
rect 60 -195 100 -185
rect 60 -265 70 -195
rect 90 -265 100 -195
rect 60 -275 100 -265
rect 125 -195 165 -185
rect 125 -265 135 -195
rect 155 -265 165 -195
rect 125 -275 165 -265
rect 190 -195 230 -185
rect 190 -265 200 -195
rect 220 -265 230 -195
rect 190 -275 230 -265
rect 15 -315 80 -295
rect 40 -335 80 -315
<< end >>
